module DLY4X1M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKAND2X6M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX8M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX40M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX32M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKBUFX40M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKBUFX24M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX16M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKBUFX12M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX24M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX24M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKBUFX20M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX8M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module TIEHIM (
	Y, 
	VDD, 
	VSS);
   output Y;
   inout VDD;
   inout VSS;
endmodule

module TIELOM (
	Y, 
	VDD, 
	VSS);
   output Y;
   inout VDD;
   inout VSS;
endmodule

module INVX2M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI21BX4M (
	Y, 
	B0N, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0N;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NAND3BX2M (
	Y, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module NAND2BX2M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module NOR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKNAND2X4M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND2X4M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module XNOR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI21X2M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module MXI2X1M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKNAND2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND3BX2M (
	Y, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module NAND2BX1M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module NAND3X2M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKNAND2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND3X1M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI21X2M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module CLKXOR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI2B1X1M (
	Y, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI2BB1X2M (
	Y, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module NAND2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI2B1X2M (
	Y, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI21X2M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AND2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI221XLM (
	Y, 
	C0, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NAND2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND3X4M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND3X4M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR3X4M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI21X4M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module XOR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND3BX4M (
	Y, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module INVX2M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MXI2X3M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI2BB2X1M (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module OAI21X2M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NOR2BX2M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX2M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR2X6M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX4M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX6M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX10M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX4M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX2M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKBUFX8M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module DLY1X4M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module INVXLM (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX2M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MX2X6M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MX2X2M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKMX2X6M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MX2X8M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module SDFFRQX2M (
	SI, 
	SE, 
	RN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module SDFFRQX4M (
	SI, 
	SE, 
	RN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module SDFFSQX2M (
	SN, 
	SI, 
	SE, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SN;
   input SI;
   input SE;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module NOR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module INVX4M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AND2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR2BX2M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module AO22X1M (
	Y, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module MX4X1M (
	Y, 
	S1, 
	S0, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S1;
   input S0;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AO21XLM (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module SDFFRHQX4M (
	SI, 
	SE, 
	RN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module SDFFRQX1M (
	SI, 
	SE, 
	RN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module SDFFRHQX2M (
	SI, 
	SE, 
	RN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module SDFFRHQX1M (
	SI, 
	SE, 
	RN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module SDFFRHQX8M (
	SI, 
	SE, 
	RN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module NAND3BX1M (
	Y, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module OAI2B2X1M (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NAND2BXLM (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module AOI2BB1XLM (
	Y, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module XOR2XLM (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR2BXLM (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module CLKMX2X2M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI211XLM (
	Y, 
	C0, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OA21X2M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI22X1M (
	Y, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NOR3X2M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MXI2X1M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR4BX1M (
	Y, 
	D, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module AOI31X2M (
	Y, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AND3X2M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI222X1M (
	Y, 
	C1, 
	C0, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C1;
   input C0;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND4BX1M (
	Y, 
	D, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module AO22XLM (
	Y, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI211X2M (
	Y, 
	C0, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI31X1M (
	Y, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OA22X2M (
	Y, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NAND3X2M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND2XLM (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MX2X1M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI2B11X2M (
	Y, 
	C0, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NAND2BX2M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module AOI2B1X1M (
	Y, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI221XLM (
	Y, 
	C0, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI22XLM (
	Y, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NOR2XLM (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OR2X1M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MXI2XLM (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AND2X1M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI32XLM (
	Y, 
	B1, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI222XLM (
	Y, 
	C1, 
	C0, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C1;
   input C0;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI31XLM (
	Y, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NOR2X1M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module ADDFX2M (
	S, 
	CO, 
	CI, 
	B, 
	A, 
	VDD, 
	VSS);
   output S;
   output CO;
   input CI;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX1M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKXOR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI21BX2M (
	Y, 
	B0N, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0N;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module XNOR2X1M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI21X1M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module XOR3XLM (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI21BX1M (
	Y, 
	B0N, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0N;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OA21X1M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI2BB1X1M (
	Y, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module ADDFHX4M (
	S, 
	CO, 
	CI, 
	B, 
	A, 
	VDD, 
	VSS);
   output S;
   output CO;
   input CI;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module ADDFHX2M (
	S, 
	CO, 
	CI, 
	B, 
	A, 
	VDD, 
	VSS);
   output S;
   output CO;
   input CI;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MX2XLM (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MXI2X2M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKMX2X4M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MXI2X6M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR2BX8M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module MXI2X3M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX6M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX4M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR3BX4M (
	Y, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module INVX8M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module XOR2X1M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR2X4M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND2X1M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MX2X2M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MXI2X4M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AND4X2M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI221X1M (
	Y, 
	C0, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI22X1M (
	Y, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AO2B2X2M (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NOR4X1M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI2BB1X2M (
	Y, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module NAND4X2M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR2BX1M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module AND4X1M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module SDFFQX2M (
	SI, 
	SE, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module SDFFQX1M (
	SI, 
	SE, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module SDFFRX1M (
	SI, 
	SE, 
	RN, 
	QN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output QN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module SDFFSQX1M (
	SN, 
	SI, 
	SE, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SN;
   input SI;
   input SE;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module OR3X2M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI32X1M (
	Y, 
	B1, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI33X2M (
	Y, 
	B2, 
	B1, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B2;
   input B1;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI33X2M (
	Y, 
	B2, 
	B1, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B2;
   input B1;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module ADDHX1M (
	S, 
	CO, 
	B, 
	A, 
	VDD, 
	VSS);
   output S;
   output CO;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR3X1M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND4X1M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI2BB1X1M (
	Y, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module NAND4BBX1M (
	Y, 
	D, 
	C, 
	BN, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input BN;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module AOI21X1M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI222X1M (
	Y, 
	C1, 
	C0, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C1;
   input C0;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NAND3XLM (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND4XLM (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI21XLM (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NOR4XLM (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI211X2M (
	Y, 
	C0, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI21BXLM (
	Y, 
	B0N, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0N;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NOR3BX2M (
	Y, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module AOI211X1M (
	Y, 
	C0, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX12M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI32XLM (
	Y, 
	B1, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI2BB1X2M (
	Y, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module AOI32X1M (
	Y, 
	B1, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module TLATNCAX16M (
	ECK, 
	E, 
	CK, 
	VDD, 
	VSS);
   output ECK;
   input E;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module OR4X1M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

/////////////////////////////////////////////////////////////
// Created by: Synopsys DC Expert(TM) in wire load mode
// Version   : K-2015.06
// Date      : Fri Oct  6 14:43:46 2023
/////////////////////////////////////////////////////////////
module mux2X1_1 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N0;

   assign N0 = SEL ;

   // Module instantiations
   MX2X6M U1 (
	.Y(OUT),
	.S0(N0),
	.B(IN_1),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux2X1_5 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N0;

   assign N0 = SEL ;

   // Module instantiations
   MX2X2M U1 (
	.Y(OUT),
	.S0(N0),
	.B(IN_1),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux2X1_4 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N0;

   assign N0 = SEL ;

   // Module instantiations
   MX2X2M U1 (
	.Y(OUT),
	.S0(N0),
	.B(IN_1),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux2X1_3 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N0;

   assign N0 = SEL ;

   // Module instantiations
   MX2X2M U1 (
	.Y(OUT),
	.S0(N0),
	.B(IN_1),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux2X1_2 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN15_RST;
   wire FE_PHN14_RST;
   wire FE_PHN3_scan_rst;
   wire FE_PHN0_scan_rst;
   wire N0;

   assign N0 = SEL ;

   // Module instantiations
   DLY4X1M FE_PHC15_RST (
	.Y(FE_PHN15_RST),
	.A(FE_PHN14_RST), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC14_RST (
	.Y(FE_PHN14_RST),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC3_scan_rst (
	.Y(FE_PHN3_scan_rst),
	.A(FE_PHN0_scan_rst), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC0_scan_rst (
	.Y(FE_PHN0_scan_rst),
	.A(IN_1), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U1 (
	.Y(OUT),
	.S0(N0),
	.B(FE_PHN3_scan_rst),
	.A(FE_PHN15_RST), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux2X1_0 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN5_scan_rst;
   wire FE_PHN2_scan_rst;
   wire N0;

   assign N0 = SEL ;

   // Module instantiations
   DLY4X1M FE_PHC5_scan_rst (
	.Y(FE_PHN5_scan_rst),
	.A(FE_PHN2_scan_rst), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC2_scan_rst (
	.Y(FE_PHN2_scan_rst),
	.A(IN_1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X6M U1 (
	.Y(OUT),
	.S0(N0),
	.B(FE_PHN5_scan_rst),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux2X1_6 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN4_scan_rst;
   wire FE_PHN1_scan_rst;
   wire N0;

   assign N0 = SEL ;

   // Module instantiations
   DLY4X1M FE_PHC4_scan_rst (
	.Y(FE_PHN4_scan_rst),
	.A(FE_PHN1_scan_rst), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC1_scan_rst (
	.Y(FE_PHN1_scan_rst),
	.A(IN_1), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X8M U1 (
	.Y(OUT),
	.S0(N0),
	.B(FE_PHN4_scan_rst),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module RegisterFile_test_1 (
	WrData, 
	Address, 
	WrEn, 
	RdEn, 
	CLK, 
	RST, 
	RdData, 
	RdData_Valid, 
	REG0, 
	REG1, 
	REG2, 
	REG3, 
	test_si2, 
	test_si1, 
	test_so2, 
	test_so1, 
	test_se, 
	FE_OFN0_rst_from_sync1, 
	FE_OFN1_rst_from_sync1, 
	ref_clock__L5_N4, 
	ref_clock__L5_N5, 
	ref_clock__L5_N6, 
	ref_clock__L5_N7, 
	VDD, 
	VSS);
   input [7:0] WrData;
   input [3:0] Address;
   input WrEn;
   input RdEn;
   input CLK;
   input RST;
   output [7:0] RdData;
   output RdData_Valid;
   output [7:0] REG0;
   output [7:0] REG1;
   output [7:0] REG2;
   output [7:0] REG3;
   input test_si2;
   input test_si1;
   output test_so2;
   output test_so1;
   input test_se;
   input FE_OFN0_rst_from_sync1;
   input FE_OFN1_rst_from_sync1;
   input ref_clock__L5_N4;
   input ref_clock__L5_N5;
   input ref_clock__L5_N6;
   input ref_clock__L5_N7;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN11_SI_2_;
   wire FE_PHN10_SI_2_;
   wire N11;
   wire N12;
   wire N13;
   wire N14;
   wire \mem[15][7] ;
   wire \mem[15][6] ;
   wire \mem[15][5] ;
   wire \mem[15][4] ;
   wire \mem[15][3] ;
   wire \mem[15][2] ;
   wire \mem[15][1] ;
   wire \mem[15][0] ;
   wire \mem[14][7] ;
   wire \mem[14][6] ;
   wire \mem[14][5] ;
   wire \mem[14][4] ;
   wire \mem[14][3] ;
   wire \mem[14][2] ;
   wire \mem[14][1] ;
   wire \mem[14][0] ;
   wire \mem[13][7] ;
   wire \mem[13][6] ;
   wire \mem[13][5] ;
   wire \mem[13][4] ;
   wire \mem[13][3] ;
   wire \mem[13][2] ;
   wire \mem[13][1] ;
   wire \mem[13][0] ;
   wire \mem[12][7] ;
   wire \mem[12][6] ;
   wire \mem[12][5] ;
   wire \mem[12][4] ;
   wire \mem[12][3] ;
   wire \mem[12][2] ;
   wire \mem[12][1] ;
   wire \mem[12][0] ;
   wire \mem[11][7] ;
   wire \mem[11][6] ;
   wire \mem[11][5] ;
   wire \mem[11][4] ;
   wire \mem[11][3] ;
   wire \mem[11][2] ;
   wire \mem[11][1] ;
   wire \mem[11][0] ;
   wire \mem[10][7] ;
   wire \mem[10][6] ;
   wire \mem[10][5] ;
   wire \mem[10][4] ;
   wire \mem[10][3] ;
   wire \mem[10][2] ;
   wire \mem[10][1] ;
   wire \mem[10][0] ;
   wire \mem[9][7] ;
   wire \mem[9][6] ;
   wire \mem[9][5] ;
   wire \mem[9][4] ;
   wire \mem[9][3] ;
   wire \mem[9][2] ;
   wire \mem[9][1] ;
   wire \mem[9][0] ;
   wire \mem[8][7] ;
   wire \mem[8][6] ;
   wire \mem[8][5] ;
   wire \mem[8][4] ;
   wire \mem[8][3] ;
   wire \mem[8][2] ;
   wire \mem[8][1] ;
   wire \mem[8][0] ;
   wire \mem[7][7] ;
   wire \mem[7][6] ;
   wire \mem[7][5] ;
   wire \mem[7][4] ;
   wire \mem[7][3] ;
   wire \mem[7][2] ;
   wire \mem[7][1] ;
   wire \mem[7][0] ;
   wire \mem[6][7] ;
   wire \mem[6][6] ;
   wire \mem[6][5] ;
   wire \mem[6][4] ;
   wire \mem[6][3] ;
   wire \mem[6][2] ;
   wire \mem[6][1] ;
   wire \mem[6][0] ;
   wire \mem[5][7] ;
   wire \mem[5][6] ;
   wire \mem[5][5] ;
   wire \mem[5][4] ;
   wire \mem[5][3] ;
   wire \mem[5][2] ;
   wire \mem[5][1] ;
   wire \mem[5][0] ;
   wire \mem[4][7] ;
   wire \mem[4][6] ;
   wire \mem[4][5] ;
   wire \mem[4][4] ;
   wire \mem[4][3] ;
   wire \mem[4][2] ;
   wire \mem[4][1] ;
   wire \mem[4][0] ;
   wire N36;
   wire N37;
   wire N38;
   wire N39;
   wire N40;
   wire N41;
   wire N42;
   wire N43;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n161;
   wire n162;
   wire n163;
   wire n164;
   wire n165;
   wire n166;
   wire n167;
   wire n168;
   wire n169;
   wire n170;
   wire n171;
   wire n172;
   wire n173;
   wire n174;
   wire n175;
   wire n176;
   wire n177;
   wire n178;
   wire n179;
   wire n180;
   wire n181;
   wire n182;
   wire n183;
   wire n184;
   wire n185;
   wire n186;
   wire n187;
   wire n188;
   wire n189;
   wire n190;
   wire n191;
   wire n192;
   wire n193;
   wire n194;
   wire n195;
   wire n196;
   wire n197;
   wire n198;
   wire n199;
   wire n200;
   wire n201;
   wire n202;
   wire n203;
   wire n204;
   wire n205;
   wire n206;
   wire n207;
   wire n208;
   wire n209;
   wire n210;
   wire n211;
   wire n212;
   wire n213;
   wire n214;
   wire n215;
   wire n216;
   wire n217;
   wire n218;
   wire n219;
   wire n220;
   wire n221;
   wire n222;
   wire n223;
   wire n224;
   wire n225;
   wire n226;
   wire n227;
   wire n228;
   wire n229;
   wire n230;
   wire n231;
   wire n232;
   wire n233;
   wire n234;
   wire n235;
   wire n236;
   wire n237;
   wire n238;
   wire n239;
   wire n240;
   wire n241;
   wire n242;
   wire n243;
   wire n244;
   wire n245;
   wire n246;
   wire n247;
   wire n248;
   wire n249;
   wire n250;
   wire n251;
   wire n252;
   wire n253;
   wire n254;
   wire n255;
   wire n256;
   wire n257;
   wire n258;
   wire n259;
   wire n260;
   wire n261;
   wire n262;
   wire n263;
   wire n264;
   wire n265;
   wire n266;
   wire n267;
   wire n268;
   wire n269;
   wire n270;
   wire n271;
   wire n272;
   wire n273;
   wire n274;
   wire n275;
   wire n276;
   wire n277;
   wire n278;
   wire n279;
   wire n280;
   wire n281;
   wire n282;
   wire n283;
   wire n284;
   wire n285;
   wire n286;
   wire n287;
   wire n288;
   wire n289;
   wire n290;
   wire n291;
   wire n292;
   wire n293;
   wire n294;
   wire n295;
   wire n296;
   wire n297;
   wire n298;
   wire n299;
   wire n300;
   wire n301;
   wire n302;
   wire n303;
   wire n304;
   wire n305;
   wire n306;
   wire n307;
   wire n308;
   wire n309;
   wire n310;
   wire n311;
   wire n312;
   wire n313;
   wire n314;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n315;
   wire n316;
   wire n317;
   wire n318;
   wire n319;
   wire n320;
   wire n321;
   wire n322;
   wire n323;
   wire n324;
   wire n325;
   wire n326;
   wire n327;
   wire n328;
   wire n329;
   wire n330;
   wire n331;
   wire n332;
   wire n333;
   wire n334;
   wire n336;
   wire n338;
   wire n339;
   wire n340;
   wire n341;
   wire n357;
   wire n358;
   wire n359;
   wire n360;
   wire n361;
   wire n362;
   wire n363;
   wire n364;
   wire n365;
   wire n366;
   wire n370;
   wire n371;
   wire n372;
   wire n373;

   assign N11 = Address[0] ;
   assign N12 = Address[1] ;
   assign N13 = Address[2] ;
   assign N14 = Address[3] ;
   assign test_so2 = \mem[15][7]  ;
   assign test_so1 = \mem[9][3]  ;

   // Module instantiations
   DLY4X1M FE_PHC11_SI_2_ (
	.Y(FE_PHN11_SI_2_),
	.A(FE_PHN10_SI_2_), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC10_SI_2_ (
	.Y(FE_PHN10_SI_2_),
	.A(test_si2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[0][7]  (
	.SI(REG0[6]),
	.SE(n370),
	.RN(RST),
	.Q(REG0[7]),
	.D(n194),
	.CK(ref_clock__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[1][0]  (
	.SI(REG0[7]),
	.SE(n373),
	.RN(RST),
	.Q(REG1[0]),
	.D(n195),
	.CK(ref_clock__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[1][7]  (
	.SI(REG1[6]),
	.SE(n372),
	.RN(RST),
	.Q(REG1[7]),
	.D(n202),
	.CK(ref_clock__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RdData_reg[0]  (
	.SI(RdData_Valid),
	.SE(n371),
	.RN(FE_OFN1_rst_from_sync1),
	.Q(RdData[0]),
	.D(n179),
	.CK(ref_clock__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[13][7]  (
	.SI(\mem[13][6] ),
	.SE(n370),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[13][7] ),
	.D(n298),
	.CK(ref_clock__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[13][6]  (
	.SI(\mem[13][5] ),
	.SE(n373),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[13][6] ),
	.D(n297),
	.CK(ref_clock__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[13][5]  (
	.SI(\mem[13][4] ),
	.SE(n372),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[13][5] ),
	.D(n296),
	.CK(ref_clock__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[13][4]  (
	.SI(\mem[13][3] ),
	.SE(n371),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[13][4] ),
	.D(n295),
	.CK(ref_clock__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[13][3]  (
	.SI(\mem[13][2] ),
	.SE(n370),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[13][3] ),
	.D(n294),
	.CK(ref_clock__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[13][2]  (
	.SI(\mem[13][1] ),
	.SE(n373),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[13][2] ),
	.D(n293),
	.CK(ref_clock__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[13][1]  (
	.SI(\mem[13][0] ),
	.SE(n372),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[13][1] ),
	.D(n292),
	.CK(ref_clock__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[13][0]  (
	.SI(\mem[12][7] ),
	.SE(n371),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[13][0] ),
	.D(n291),
	.CK(ref_clock__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[9][7]  (
	.SI(\mem[9][6] ),
	.SE(n370),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[9][7] ),
	.D(n266),
	.CK(ref_clock__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[9][6]  (
	.SI(\mem[9][5] ),
	.SE(n373),
	.RN(FE_OFN1_rst_from_sync1),
	.Q(\mem[9][6] ),
	.D(n265),
	.CK(ref_clock__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[9][5]  (
	.SI(\mem[9][4] ),
	.SE(n372),
	.RN(FE_OFN1_rst_from_sync1),
	.Q(\mem[9][5] ),
	.D(n264),
	.CK(ref_clock__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[9][4]  (
	.SI(FE_PHN11_SI_2_),
	.SE(n371),
	.RN(FE_OFN1_rst_from_sync1),
	.Q(\mem[9][4] ),
	.D(n263),
	.CK(ref_clock__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX4M \mem_reg[9][3]  (
	.SI(\mem[9][2] ),
	.SE(n370),
	.RN(FE_OFN1_rst_from_sync1),
	.Q(\mem[9][3] ),
	.D(n262),
	.CK(ref_clock__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[9][2]  (
	.SI(\mem[9][1] ),
	.SE(n373),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[9][2] ),
	.D(n261),
	.CK(ref_clock__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[9][1]  (
	.SI(\mem[9][0] ),
	.SE(n372),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[9][1] ),
	.D(n260),
	.CK(ref_clock__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[9][0]  (
	.SI(\mem[8][7] ),
	.SE(n371),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[9][0] ),
	.D(n259),
	.CK(ref_clock__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[5][7]  (
	.SI(\mem[5][6] ),
	.SE(n370),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[5][7] ),
	.D(n234),
	.CK(ref_clock__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[5][6]  (
	.SI(\mem[5][5] ),
	.SE(n373),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[5][6] ),
	.D(n233),
	.CK(ref_clock__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[5][5]  (
	.SI(\mem[5][4] ),
	.SE(n372),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[5][5] ),
	.D(n232),
	.CK(ref_clock__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[5][4]  (
	.SI(\mem[5][3] ),
	.SE(n371),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[5][4] ),
	.D(n231),
	.CK(ref_clock__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[5][3]  (
	.SI(\mem[5][2] ),
	.SE(n370),
	.RN(RST),
	.Q(\mem[5][3] ),
	.D(n230),
	.CK(ref_clock__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[5][2]  (
	.SI(\mem[5][1] ),
	.SE(n373),
	.RN(RST),
	.Q(\mem[5][2] ),
	.D(n229),
	.CK(ref_clock__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[5][1]  (
	.SI(\mem[5][0] ),
	.SE(n372),
	.RN(RST),
	.Q(\mem[5][1] ),
	.D(n228),
	.CK(ref_clock__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[5][0]  (
	.SI(\mem[4][7] ),
	.SE(n371),
	.RN(RST),
	.Q(\mem[5][0] ),
	.D(n227),
	.CK(ref_clock__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[15][7]  (
	.SI(\mem[15][6] ),
	.SE(n370),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[15][7] ),
	.D(n314),
	.CK(ref_clock__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[15][6]  (
	.SI(\mem[15][5] ),
	.SE(n373),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[15][6] ),
	.D(n313),
	.CK(ref_clock__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[15][5]  (
	.SI(\mem[15][4] ),
	.SE(n372),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[15][5] ),
	.D(n312),
	.CK(ref_clock__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[15][4]  (
	.SI(\mem[15][3] ),
	.SE(n371),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[15][4] ),
	.D(n311),
	.CK(ref_clock__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[15][3]  (
	.SI(\mem[15][2] ),
	.SE(n370),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[15][3] ),
	.D(n310),
	.CK(ref_clock__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[15][2]  (
	.SI(\mem[15][1] ),
	.SE(n373),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[15][2] ),
	.D(n309),
	.CK(ref_clock__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[15][1]  (
	.SI(\mem[15][0] ),
	.SE(n372),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[15][1] ),
	.D(n308),
	.CK(ref_clock__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[15][0]  (
	.SI(\mem[14][7] ),
	.SE(n371),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[15][0] ),
	.D(n307),
	.CK(ref_clock__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[11][7]  (
	.SI(\mem[11][6] ),
	.SE(n370),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[11][7] ),
	.D(n282),
	.CK(ref_clock__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[11][6]  (
	.SI(\mem[11][5] ),
	.SE(n373),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[11][6] ),
	.D(n281),
	.CK(ref_clock__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[11][5]  (
	.SI(\mem[11][4] ),
	.SE(n372),
	.RN(FE_OFN1_rst_from_sync1),
	.Q(\mem[11][5] ),
	.D(n280),
	.CK(ref_clock__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[11][4]  (
	.SI(\mem[11][3] ),
	.SE(n371),
	.RN(FE_OFN1_rst_from_sync1),
	.Q(\mem[11][4] ),
	.D(n279),
	.CK(ref_clock__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[11][3]  (
	.SI(\mem[11][2] ),
	.SE(n370),
	.RN(FE_OFN1_rst_from_sync1),
	.Q(\mem[11][3] ),
	.D(n278),
	.CK(ref_clock__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[11][2]  (
	.SI(\mem[11][1] ),
	.SE(n373),
	.RN(FE_OFN1_rst_from_sync1),
	.Q(\mem[11][2] ),
	.D(n277),
	.CK(ref_clock__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[11][1]  (
	.SI(\mem[11][0] ),
	.SE(n372),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[11][1] ),
	.D(n276),
	.CK(ref_clock__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[11][0]  (
	.SI(\mem[10][7] ),
	.SE(n371),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[11][0] ),
	.D(n275),
	.CK(ref_clock__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[7][7]  (
	.SI(\mem[7][6] ),
	.SE(n370),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[7][7] ),
	.D(n250),
	.CK(ref_clock__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[7][6]  (
	.SI(\mem[7][5] ),
	.SE(n373),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[7][6] ),
	.D(n249),
	.CK(ref_clock__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[7][5]  (
	.SI(\mem[7][4] ),
	.SE(n372),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[7][5] ),
	.D(n248),
	.CK(ref_clock__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[7][4]  (
	.SI(\mem[7][3] ),
	.SE(n371),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[7][4] ),
	.D(n247),
	.CK(ref_clock__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[7][3]  (
	.SI(\mem[7][2] ),
	.SE(n370),
	.RN(RST),
	.Q(\mem[7][3] ),
	.D(n246),
	.CK(ref_clock__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[7][2]  (
	.SI(\mem[7][1] ),
	.SE(n373),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[7][2] ),
	.D(n245),
	.CK(ref_clock__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[7][1]  (
	.SI(\mem[7][0] ),
	.SE(n372),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[7][1] ),
	.D(n244),
	.CK(ref_clock__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[7][0]  (
	.SI(\mem[6][7] ),
	.SE(n371),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[7][0] ),
	.D(n243),
	.CK(ref_clock__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[14][7]  (
	.SI(\mem[14][6] ),
	.SE(n370),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[14][7] ),
	.D(n306),
	.CK(ref_clock__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[14][6]  (
	.SI(\mem[14][5] ),
	.SE(n373),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[14][6] ),
	.D(n305),
	.CK(ref_clock__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[14][5]  (
	.SI(\mem[14][4] ),
	.SE(n372),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[14][5] ),
	.D(n304),
	.CK(ref_clock__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[14][4]  (
	.SI(\mem[14][3] ),
	.SE(n371),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[14][4] ),
	.D(n303),
	.CK(ref_clock__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[14][3]  (
	.SI(\mem[14][2] ),
	.SE(n370),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[14][3] ),
	.D(n302),
	.CK(ref_clock__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[14][2]  (
	.SI(\mem[14][1] ),
	.SE(n373),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[14][2] ),
	.D(n301),
	.CK(ref_clock__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[14][1]  (
	.SI(\mem[14][0] ),
	.SE(n372),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[14][1] ),
	.D(n300),
	.CK(ref_clock__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[14][0]  (
	.SI(\mem[13][7] ),
	.SE(n371),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[14][0] ),
	.D(n299),
	.CK(ref_clock__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[10][7]  (
	.SI(\mem[10][6] ),
	.SE(n370),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[10][7] ),
	.D(n274),
	.CK(ref_clock__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[10][6]  (
	.SI(\mem[10][5] ),
	.SE(n373),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[10][6] ),
	.D(n273),
	.CK(ref_clock__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[10][5]  (
	.SI(\mem[10][4] ),
	.SE(n372),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[10][5] ),
	.D(n272),
	.CK(ref_clock__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[10][4]  (
	.SI(\mem[10][3] ),
	.SE(n371),
	.RN(FE_OFN1_rst_from_sync1),
	.Q(\mem[10][4] ),
	.D(n271),
	.CK(ref_clock__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[10][3]  (
	.SI(\mem[10][2] ),
	.SE(n370),
	.RN(FE_OFN1_rst_from_sync1),
	.Q(\mem[10][3] ),
	.D(n270),
	.CK(ref_clock__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[10][2]  (
	.SI(\mem[10][1] ),
	.SE(n373),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[10][2] ),
	.D(n269),
	.CK(ref_clock__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[10][1]  (
	.SI(\mem[10][0] ),
	.SE(n372),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[10][1] ),
	.D(n268),
	.CK(ref_clock__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[10][0]  (
	.SI(\mem[9][7] ),
	.SE(n371),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[10][0] ),
	.D(n267),
	.CK(ref_clock__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[6][7]  (
	.SI(\mem[6][6] ),
	.SE(n370),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[6][7] ),
	.D(n242),
	.CK(ref_clock__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[6][6]  (
	.SI(\mem[6][5] ),
	.SE(n373),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[6][6] ),
	.D(n241),
	.CK(ref_clock__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[6][5]  (
	.SI(\mem[6][4] ),
	.SE(n372),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[6][5] ),
	.D(n240),
	.CK(ref_clock__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[6][4]  (
	.SI(\mem[6][3] ),
	.SE(n371),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[6][4] ),
	.D(n239),
	.CK(ref_clock__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[6][3]  (
	.SI(\mem[6][2] ),
	.SE(n370),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[6][3] ),
	.D(n238),
	.CK(ref_clock__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[6][2]  (
	.SI(\mem[6][1] ),
	.SE(n373),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[6][2] ),
	.D(n237),
	.CK(ref_clock__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[6][1]  (
	.SI(\mem[6][0] ),
	.SE(n372),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[6][1] ),
	.D(n236),
	.CK(ref_clock__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[6][0]  (
	.SI(\mem[5][7] ),
	.SE(n371),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[6][0] ),
	.D(n235),
	.CK(ref_clock__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[12][7]  (
	.SI(\mem[12][6] ),
	.SE(n370),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[12][7] ),
	.D(n290),
	.CK(ref_clock__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[12][6]  (
	.SI(\mem[12][5] ),
	.SE(n373),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[12][6] ),
	.D(n289),
	.CK(ref_clock__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[12][5]  (
	.SI(\mem[12][4] ),
	.SE(n372),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[12][5] ),
	.D(n288),
	.CK(ref_clock__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[12][4]  (
	.SI(\mem[12][3] ),
	.SE(n371),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[12][4] ),
	.D(n287),
	.CK(ref_clock__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[12][3]  (
	.SI(\mem[12][2] ),
	.SE(n370),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[12][3] ),
	.D(n286),
	.CK(ref_clock__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[12][2]  (
	.SI(\mem[12][1] ),
	.SE(n373),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[12][2] ),
	.D(n285),
	.CK(ref_clock__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[12][1]  (
	.SI(\mem[12][0] ),
	.SE(n372),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[12][1] ),
	.D(n284),
	.CK(ref_clock__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[12][0]  (
	.SI(\mem[11][7] ),
	.SE(n371),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[12][0] ),
	.D(n283),
	.CK(ref_clock__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[8][7]  (
	.SI(\mem[8][6] ),
	.SE(n370),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[8][7] ),
	.D(n258),
	.CK(ref_clock__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[8][6]  (
	.SI(\mem[8][5] ),
	.SE(n373),
	.RN(FE_OFN1_rst_from_sync1),
	.Q(\mem[8][6] ),
	.D(n257),
	.CK(ref_clock__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[8][5]  (
	.SI(\mem[8][4] ),
	.SE(n372),
	.RN(FE_OFN1_rst_from_sync1),
	.Q(\mem[8][5] ),
	.D(n256),
	.CK(ref_clock__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[8][4]  (
	.SI(\mem[8][3] ),
	.SE(n371),
	.RN(FE_OFN1_rst_from_sync1),
	.Q(\mem[8][4] ),
	.D(n255),
	.CK(ref_clock__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[8][3]  (
	.SI(\mem[8][2] ),
	.SE(n370),
	.RN(FE_OFN1_rst_from_sync1),
	.Q(\mem[8][3] ),
	.D(n254),
	.CK(ref_clock__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[8][2]  (
	.SI(\mem[8][1] ),
	.SE(n373),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[8][2] ),
	.D(n253),
	.CK(ref_clock__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[8][1]  (
	.SI(\mem[8][0] ),
	.SE(n372),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[8][1] ),
	.D(n252),
	.CK(ref_clock__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[8][0]  (
	.SI(\mem[7][7] ),
	.SE(n371),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[8][0] ),
	.D(n251),
	.CK(ref_clock__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[4][7]  (
	.SI(\mem[4][6] ),
	.SE(n370),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[4][7] ),
	.D(n226),
	.CK(ref_clock__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[4][6]  (
	.SI(\mem[4][5] ),
	.SE(n373),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[4][6] ),
	.D(n225),
	.CK(ref_clock__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[4][5]  (
	.SI(\mem[4][4] ),
	.SE(n372),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[4][5] ),
	.D(n224),
	.CK(ref_clock__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[4][4]  (
	.SI(\mem[4][3] ),
	.SE(n371),
	.RN(FE_OFN0_rst_from_sync1),
	.Q(\mem[4][4] ),
	.D(n223),
	.CK(ref_clock__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[4][3]  (
	.SI(\mem[4][2] ),
	.SE(n370),
	.RN(RST),
	.Q(\mem[4][3] ),
	.D(n222),
	.CK(ref_clock__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[4][2]  (
	.SI(\mem[4][1] ),
	.SE(n373),
	.RN(RST),
	.Q(\mem[4][2] ),
	.D(n221),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[4][1]  (
	.SI(\mem[4][0] ),
	.SE(n372),
	.RN(RST),
	.Q(\mem[4][1] ),
	.D(n220),
	.CK(ref_clock__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[4][0]  (
	.SI(REG3[7]),
	.SE(n371),
	.RN(RST),
	.Q(\mem[4][0] ),
	.D(n219),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[1][5]  (
	.SI(REG1[4]),
	.SE(n370),
	.RN(FE_OFN1_rst_from_sync1),
	.Q(REG1[5]),
	.D(n200),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[1][4]  (
	.SI(REG1[3]),
	.SE(n373),
	.RN(FE_OFN1_rst_from_sync1),
	.Q(REG1[4]),
	.D(n199),
	.CK(ref_clock__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[1][3]  (
	.SI(REG1[2]),
	.SE(n372),
	.RN(FE_OFN1_rst_from_sync1),
	.Q(REG1[3]),
	.D(n198),
	.CK(ref_clock__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[1][2]  (
	.SI(REG1[1]),
	.SE(n371),
	.RN(FE_OFN1_rst_from_sync1),
	.Q(REG1[2]),
	.D(n197),
	.CK(ref_clock__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[1][1]  (
	.SI(REG1[0]),
	.SE(n370),
	.RN(FE_OFN1_rst_from_sync1),
	.Q(REG1[1]),
	.D(n196),
	.CK(ref_clock__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[1][6]  (
	.SI(REG1[5]),
	.SE(n373),
	.RN(RST),
	.Q(REG1[6]),
	.D(n201),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[0][6]  (
	.SI(REG0[5]),
	.SE(n372),
	.RN(FE_OFN1_rst_from_sync1),
	.Q(REG0[6]),
	.D(n193),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[0][5]  (
	.SI(REG0[4]),
	.SE(n371),
	.RN(FE_OFN1_rst_from_sync1),
	.Q(REG0[5]),
	.D(n192),
	.CK(ref_clock__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[0][4]  (
	.SI(REG0[3]),
	.SE(n370),
	.RN(FE_OFN1_rst_from_sync1),
	.Q(REG0[4]),
	.D(n191),
	.CK(ref_clock__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[0][3]  (
	.SI(REG0[2]),
	.SE(n373),
	.RN(FE_OFN1_rst_from_sync1),
	.Q(REG0[3]),
	.D(n190),
	.CK(ref_clock__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[0][2]  (
	.SI(REG0[1]),
	.SE(n372),
	.RN(FE_OFN1_rst_from_sync1),
	.Q(REG0[2]),
	.D(n189),
	.CK(ref_clock__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[0][1]  (
	.SI(REG0[0]),
	.SE(n371),
	.RN(FE_OFN1_rst_from_sync1),
	.Q(REG0[1]),
	.D(n188),
	.CK(ref_clock__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[0][0]  (
	.SI(RdData[7]),
	.SE(n370),
	.RN(FE_OFN1_rst_from_sync1),
	.Q(REG0[0]),
	.D(n187),
	.CK(ref_clock__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RdData_reg[7]  (
	.SI(RdData[6]),
	.SE(n373),
	.RN(FE_OFN1_rst_from_sync1),
	.Q(RdData[7]),
	.D(n186),
	.CK(ref_clock__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RdData_reg[6]  (
	.SI(RdData[5]),
	.SE(n372),
	.RN(FE_OFN1_rst_from_sync1),
	.Q(RdData[6]),
	.D(n185),
	.CK(ref_clock__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RdData_reg[5]  (
	.SI(RdData[4]),
	.SE(n371),
	.RN(FE_OFN1_rst_from_sync1),
	.Q(RdData[5]),
	.D(n184),
	.CK(ref_clock__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RdData_reg[4]  (
	.SI(RdData[3]),
	.SE(n370),
	.RN(FE_OFN1_rst_from_sync1),
	.Q(RdData[4]),
	.D(n183),
	.CK(ref_clock__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RdData_reg[3]  (
	.SI(RdData[2]),
	.SE(n373),
	.RN(FE_OFN1_rst_from_sync1),
	.Q(RdData[3]),
	.D(n182),
	.CK(ref_clock__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RdData_reg[2]  (
	.SI(RdData[1]),
	.SE(n372),
	.RN(FE_OFN1_rst_from_sync1),
	.Q(RdData[2]),
	.D(n181),
	.CK(ref_clock__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RdData_reg[1]  (
	.SI(RdData[0]),
	.SE(n371),
	.RN(FE_OFN1_rst_from_sync1),
	.Q(RdData[1]),
	.D(n180),
	.CK(ref_clock__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[2][1]  (
	.SI(REG2[0]),
	.SE(n370),
	.RN(RST),
	.Q(REG2[1]),
	.D(n204),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSQX2M \mem_reg[2][0]  (
	.SN(RST),
	.SI(REG1[7]),
	.SE(n373),
	.Q(REG2[0]),
	.D(n203),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[3][0]  (
	.SI(REG2[7]),
	.SE(n373),
	.RN(RST),
	.Q(REG3[0]),
	.D(n211),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M RdData_Valid_reg (
	.SI(test_si1),
	.SE(n372),
	.RN(FE_OFN1_rst_from_sync1),
	.Q(RdData_Valid),
	.D(n178),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[3][1]  (
	.SI(REG3[0]),
	.SE(n371),
	.RN(RST),
	.Q(REG3[1]),
	.D(n212),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSQX2M \mem_reg[3][5]  (
	.SN(RST),
	.SI(REG3[4]),
	.SE(n372),
	.Q(REG3[5]),
	.D(n216),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[3][4]  (
	.SI(REG3[3]),
	.SE(n370),
	.RN(RST),
	.Q(REG3[4]),
	.D(n215),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[3][3]  (
	.SI(REG3[2]),
	.SE(n373),
	.RN(RST),
	.Q(REG3[3]),
	.D(n214),
	.CK(ref_clock__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[3][2]  (
	.SI(REG3[1]),
	.SE(n372),
	.RN(RST),
	.Q(REG3[2]),
	.D(n213),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[3][6]  (
	.SI(REG3[5]),
	.SE(n371),
	.RN(RST),
	.Q(REG3[6]),
	.D(n217),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[3][7]  (
	.SI(REG3[6]),
	.SE(n370),
	.RN(RST),
	.Q(REG3[7]),
	.D(n218),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[2][2]  (
	.SI(REG2[1]),
	.SE(n373),
	.RN(RST),
	.Q(REG2[2]),
	.D(n205),
	.CK(ref_clock__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[2][3]  (
	.SI(REG2[2]),
	.SE(n372),
	.RN(RST),
	.Q(REG2[3]),
	.D(n206),
	.CK(ref_clock__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSQX2M \mem_reg[2][7]  (
	.SN(RST),
	.SI(REG2[6]),
	.SE(n371),
	.Q(REG2[7]),
	.D(n210),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[2][4]  (
	.SI(REG2[3]),
	.SE(n371),
	.RN(RST),
	.Q(REG2[4]),
	.D(n207),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[2][6]  (
	.SI(REG2[5]),
	.SE(n370),
	.RN(RST),
	.Q(REG2[6]),
	.D(n209),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[2][5]  (
	.SI(REG2[4]),
	.SE(test_se),
	.RN(RST),
	.Q(REG2[5]),
	.D(n208),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U140 (
	.Y(n153),
	.B(N13),
	.A(N12), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U141 (
	.Y(n158),
	.B(N13),
	.A(n341), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX4M U142 (
	.Y(n338),
	.A(n340), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U143 (
	.Y(n336),
	.A(n341), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX4M U144 (
	.Y(n339),
	.A(n340), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U147 (
	.Y(n155),
	.B(n153),
	.A(n156), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U148 (
	.Y(n167),
	.B(n153),
	.A(n168), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U149 (
	.Y(n169),
	.B(n153),
	.A(n170), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U150 (
	.Y(n171),
	.B(n158),
	.A(n168), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U151 (
	.Y(n172),
	.B(n158),
	.A(n170), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U152 (
	.Y(n157),
	.B(n154),
	.A(n158), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U153 (
	.Y(n159),
	.B(n156),
	.A(n158), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U154 (
	.Y(n160),
	.B(n154),
	.A(n161), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U155 (
	.Y(n162),
	.B(n156),
	.A(n161), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U156 (
	.Y(n163),
	.B(n154),
	.A(n164), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U157 (
	.Y(n166),
	.B(n156),
	.A(n164), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U158 (
	.Y(n173),
	.B(n161),
	.A(n168), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U159 (
	.Y(n174),
	.B(n161),
	.A(n170), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U160 (
	.Y(n175),
	.B(n164),
	.A(n168), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U161 (
	.Y(n177),
	.B(n164),
	.A(n170), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U162 (
	.Y(n152),
	.B(n154),
	.A(n153), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U163 (
	.Y(n154),
	.B(n340),
	.A(n165), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U164 (
	.Y(n156),
	.B(N11),
	.A(n165), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U165 (
	.Y(n168),
	.B(n340),
	.A(n176), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U166 (
	.Y(n170),
	.B(N11),
	.A(n176), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U167 (
	.Y(n357),
	.A(n151), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U178 (
	.Y(n340),
	.A(N11), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U179 (
	.Y(n359),
	.A(WrData[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U180 (
	.Y(n360),
	.A(WrData[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U181 (
	.Y(n361),
	.A(WrData[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U182 (
	.Y(n362),
	.A(WrData[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U183 (
	.Y(n363),
	.A(WrData[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U184 (
	.Y(n364),
	.A(WrData[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U185 (
	.Y(n365),
	.A(WrData[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U186 (
	.Y(n366),
	.A(WrData[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U187 (
	.Y(n151),
	.B(n358),
	.A(RdEn), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U188 (
	.Y(n165),
	.B(N14),
	.AN(n150), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U189 (
	.Y(n150),
	.B(RdEn),
	.A(n358), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U190 (
	.Y(n161),
	.B(n341),
	.A(N13), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U191 (
	.Y(n164),
	.B(N12),
	.A(N13), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U192 (
	.Y(n176),
	.B(n150),
	.A(N14), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U193 (
	.Y(n341),
	.A(N12), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U199 (
	.Y(n179),
	.B1(n151),
	.B0(RdData[0]),
	.A1(n357),
	.A0(N43), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U200 (
	.Y(N43),
	.S1(N13),
	.S0(N14),
	.D(n138),
	.C(n140),
	.B(n139),
	.A(n141), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U201 (
	.Y(n141),
	.S1(N12),
	.S0(N11),
	.D(REG3[0]),
	.C(REG2[0]),
	.B(REG1[0]),
	.A(REG0[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U202 (
	.Y(n139),
	.S1(N12),
	.S0(N11),
	.D(\mem[11][0] ),
	.C(\mem[10][0] ),
	.B(\mem[9][0] ),
	.A(\mem[8][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U203 (
	.Y(n180),
	.B1(n151),
	.B0(RdData[1]),
	.A1(n357),
	.A0(N42), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U204 (
	.Y(N42),
	.S1(N13),
	.S0(N14),
	.D(n142),
	.C(n144),
	.B(n143),
	.A(n145), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U205 (
	.Y(n143),
	.S1(N12),
	.S0(N11),
	.D(\mem[11][1] ),
	.C(\mem[10][1] ),
	.B(\mem[9][1] ),
	.A(\mem[8][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U206 (
	.Y(n142),
	.S1(n336),
	.S0(n339),
	.D(\mem[15][1] ),
	.C(\mem[14][1] ),
	.B(\mem[13][1] ),
	.A(\mem[12][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U207 (
	.Y(n181),
	.B1(n151),
	.B0(RdData[2]),
	.A1(n357),
	.A0(N41), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U208 (
	.Y(N41),
	.S1(N13),
	.S0(N14),
	.D(n146),
	.C(n148),
	.B(n147),
	.A(n149), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U209 (
	.Y(n149),
	.S1(n336),
	.S0(n338),
	.D(REG3[2]),
	.C(REG2[2]),
	.B(REG1[2]),
	.A(REG0[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U210 (
	.Y(n147),
	.S1(n336),
	.S0(n338),
	.D(\mem[11][2] ),
	.C(\mem[10][2] ),
	.B(\mem[9][2] ),
	.A(\mem[8][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U211 (
	.Y(n182),
	.B1(n151),
	.B0(RdData[3]),
	.A1(n357),
	.A0(N40), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U212 (
	.Y(N40),
	.S1(N13),
	.S0(N14),
	.D(n315),
	.C(n317),
	.B(n316),
	.A(n318), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U213 (
	.Y(n318),
	.S1(n336),
	.S0(n338),
	.D(REG3[3]),
	.C(REG2[3]),
	.B(REG1[3]),
	.A(REG0[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U214 (
	.Y(n316),
	.S1(n336),
	.S0(n338),
	.D(\mem[11][3] ),
	.C(\mem[10][3] ),
	.B(\mem[9][3] ),
	.A(\mem[8][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U215 (
	.Y(n183),
	.B1(n151),
	.B0(RdData[4]),
	.A1(n357),
	.A0(N39), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U216 (
	.Y(N39),
	.S1(N13),
	.S0(N14),
	.D(n319),
	.C(n321),
	.B(n320),
	.A(n322), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U217 (
	.Y(n322),
	.S1(n336),
	.S0(n339),
	.D(REG3[4]),
	.C(REG2[4]),
	.B(REG1[4]),
	.A(REG0[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U218 (
	.Y(n320),
	.S1(n336),
	.S0(n338),
	.D(\mem[11][4] ),
	.C(\mem[10][4] ),
	.B(\mem[9][4] ),
	.A(\mem[8][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U219 (
	.Y(n184),
	.B1(n151),
	.B0(RdData[5]),
	.A1(n357),
	.A0(N38), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U220 (
	.Y(N38),
	.S1(N13),
	.S0(N14),
	.D(n323),
	.C(n325),
	.B(n324),
	.A(n326), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U221 (
	.Y(n326),
	.S1(N12),
	.S0(n339),
	.D(REG3[5]),
	.C(REG2[5]),
	.B(REG1[5]),
	.A(REG0[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U222 (
	.Y(n324),
	.S1(N12),
	.S0(n339),
	.D(\mem[11][5] ),
	.C(\mem[10][5] ),
	.B(\mem[9][5] ),
	.A(\mem[8][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U223 (
	.Y(n185),
	.B1(n151),
	.B0(RdData[6]),
	.A1(n357),
	.A0(N37), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U224 (
	.Y(N37),
	.S1(N13),
	.S0(N14),
	.D(n327),
	.C(n329),
	.B(n328),
	.A(n330), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U225 (
	.Y(n330),
	.S1(N12),
	.S0(n339),
	.D(REG3[6]),
	.C(REG2[6]),
	.B(REG1[6]),
	.A(REG0[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U226 (
	.Y(n328),
	.S1(N12),
	.S0(n339),
	.D(\mem[11][6] ),
	.C(\mem[10][6] ),
	.B(\mem[9][6] ),
	.A(\mem[8][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U227 (
	.Y(n186),
	.B1(n151),
	.B0(RdData[7]),
	.A1(n357),
	.A0(N36), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U228 (
	.Y(N36),
	.S1(N13),
	.S0(N14),
	.D(n331),
	.C(n333),
	.B(n332),
	.A(n334), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U229 (
	.Y(n334),
	.S1(N12),
	.S0(n339),
	.D(REG3[7]),
	.C(REG2[7]),
	.B(REG1[7]),
	.A(REG0[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U230 (
	.Y(n332),
	.S1(N12),
	.S0(n339),
	.D(\mem[11][7] ),
	.C(\mem[10][7] ),
	.B(\mem[9][7] ),
	.A(\mem[8][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U231 (
	.Y(n145),
	.S1(N12),
	.S0(n338),
	.D(REG3[1]),
	.C(REG2[1]),
	.B(REG1[1]),
	.A(REG0[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U232 (
	.Y(n140),
	.S1(N12),
	.S0(N11),
	.D(\mem[7][0] ),
	.C(\mem[6][0] ),
	.B(\mem[5][0] ),
	.A(\mem[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U233 (
	.Y(n144),
	.S1(N12),
	.S0(n338),
	.D(\mem[7][1] ),
	.C(\mem[6][1] ),
	.B(\mem[5][1] ),
	.A(\mem[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U234 (
	.Y(n148),
	.S1(n336),
	.S0(n338),
	.D(\mem[7][2] ),
	.C(\mem[6][2] ),
	.B(\mem[5][2] ),
	.A(\mem[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U235 (
	.Y(n317),
	.S1(n336),
	.S0(n338),
	.D(\mem[7][3] ),
	.C(\mem[6][3] ),
	.B(\mem[5][3] ),
	.A(\mem[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U236 (
	.Y(n321),
	.S1(n336),
	.S0(n338),
	.D(\mem[7][4] ),
	.C(\mem[6][4] ),
	.B(\mem[5][4] ),
	.A(\mem[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U237 (
	.Y(n325),
	.S1(N12),
	.S0(n339),
	.D(\mem[7][5] ),
	.C(\mem[6][5] ),
	.B(\mem[5][5] ),
	.A(\mem[4][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U238 (
	.Y(n329),
	.S1(N12),
	.S0(n339),
	.D(\mem[7][6] ),
	.C(\mem[6][6] ),
	.B(\mem[5][6] ),
	.A(\mem[4][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U239 (
	.Y(n333),
	.S1(N12),
	.S0(n339),
	.D(\mem[7][7] ),
	.C(\mem[6][7] ),
	.B(\mem[5][7] ),
	.A(\mem[4][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U240 (
	.Y(n138),
	.S1(n336),
	.S0(n338),
	.D(\mem[15][0] ),
	.C(\mem[14][0] ),
	.B(\mem[13][0] ),
	.A(\mem[12][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U241 (
	.Y(n146),
	.S1(n336),
	.S0(n338),
	.D(\mem[15][2] ),
	.C(\mem[14][2] ),
	.B(\mem[13][2] ),
	.A(\mem[12][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U242 (
	.Y(n315),
	.S1(n336),
	.S0(n338),
	.D(\mem[15][3] ),
	.C(\mem[14][3] ),
	.B(\mem[13][3] ),
	.A(\mem[12][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U243 (
	.Y(n319),
	.S1(n336),
	.S0(n338),
	.D(\mem[15][4] ),
	.C(\mem[14][4] ),
	.B(\mem[13][4] ),
	.A(\mem[12][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U244 (
	.Y(n323),
	.S1(N12),
	.S0(n339),
	.D(\mem[15][5] ),
	.C(\mem[14][5] ),
	.B(\mem[13][5] ),
	.A(\mem[12][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U245 (
	.Y(n327),
	.S1(N12),
	.S0(n339),
	.D(\mem[15][6] ),
	.C(\mem[14][6] ),
	.B(\mem[13][6] ),
	.A(\mem[12][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U246 (
	.Y(n331),
	.S1(N12),
	.S0(n339),
	.D(\mem[15][7] ),
	.C(\mem[14][7] ),
	.B(\mem[13][7] ),
	.A(\mem[12][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U247 (
	.Y(n187),
	.B1(n359),
	.B0(n152),
	.A1N(n152),
	.A0N(REG0[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U248 (
	.Y(n188),
	.B1(n360),
	.B0(n152),
	.A1N(n152),
	.A0N(REG0[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U249 (
	.Y(n189),
	.B1(n361),
	.B0(n152),
	.A1N(n152),
	.A0N(REG0[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U250 (
	.Y(n190),
	.B1(n362),
	.B0(n152),
	.A1N(n152),
	.A0N(REG0[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U251 (
	.Y(n191),
	.B1(n363),
	.B0(n152),
	.A1N(n152),
	.A0N(REG0[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U252 (
	.Y(n192),
	.B1(n364),
	.B0(n152),
	.A1N(n152),
	.A0N(REG0[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U253 (
	.Y(n193),
	.B1(n365),
	.B0(n152),
	.A1N(n152),
	.A0N(REG0[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U254 (
	.Y(n204),
	.B1(n157),
	.B0(n360),
	.A1N(n157),
	.A0N(REG2[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U255 (
	.Y(n205),
	.B1(n157),
	.B0(n361),
	.A1N(n157),
	.A0N(REG2[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U256 (
	.Y(n206),
	.B1(n157),
	.B0(n362),
	.A1N(n157),
	.A0N(REG2[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U257 (
	.Y(n207),
	.B1(n157),
	.B0(n363),
	.A1N(n157),
	.A0N(REG2[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U258 (
	.Y(n208),
	.B1(n157),
	.B0(n364),
	.A1N(n157),
	.A0N(REG2[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U259 (
	.Y(n209),
	.B1(n157),
	.B0(n365),
	.A1N(n157),
	.A0N(REG2[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U260 (
	.Y(n211),
	.B1(n159),
	.B0(n359),
	.A1N(n159),
	.A0N(REG3[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U261 (
	.Y(n212),
	.B1(n159),
	.B0(n360),
	.A1N(n159),
	.A0N(REG3[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U262 (
	.Y(n213),
	.B1(n159),
	.B0(n361),
	.A1N(n159),
	.A0N(REG3[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U263 (
	.Y(n214),
	.B1(n159),
	.B0(n362),
	.A1N(n159),
	.A0N(REG3[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U264 (
	.Y(n215),
	.B1(n159),
	.B0(n363),
	.A1N(n159),
	.A0N(REG3[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U265 (
	.Y(n217),
	.B1(n159),
	.B0(n365),
	.A1N(n159),
	.A0N(REG3[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U266 (
	.Y(n218),
	.B1(n159),
	.B0(n366),
	.A1N(n159),
	.A0N(REG3[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U267 (
	.Y(n196),
	.B1(n155),
	.B0(n360),
	.A1N(n155),
	.A0N(REG1[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U268 (
	.Y(n197),
	.B1(n155),
	.B0(n361),
	.A1N(n155),
	.A0N(REG1[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U269 (
	.Y(n198),
	.B1(n155),
	.B0(n362),
	.A1N(n155),
	.A0N(REG1[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U270 (
	.Y(n199),
	.B1(n155),
	.B0(n363),
	.A1N(n155),
	.A0N(REG1[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U271 (
	.Y(n200),
	.B1(n155),
	.B0(n364),
	.A1N(n155),
	.A0N(REG1[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U272 (
	.Y(n201),
	.B1(n155),
	.B0(n365),
	.A1N(n155),
	.A0N(REG1[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U273 (
	.Y(n251),
	.B1(n167),
	.B0(n359),
	.A1N(n167),
	.A0N(\mem[8][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U274 (
	.Y(n252),
	.B1(n167),
	.B0(n360),
	.A1N(n167),
	.A0N(\mem[8][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U275 (
	.Y(n253),
	.B1(n167),
	.B0(n361),
	.A1N(n167),
	.A0N(\mem[8][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U276 (
	.Y(n254),
	.B1(n167),
	.B0(n362),
	.A1N(n167),
	.A0N(\mem[8][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U277 (
	.Y(n255),
	.B1(n167),
	.B0(n363),
	.A1N(n167),
	.A0N(\mem[8][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U278 (
	.Y(n256),
	.B1(n167),
	.B0(n364),
	.A1N(n167),
	.A0N(\mem[8][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U279 (
	.Y(n257),
	.B1(n167),
	.B0(n365),
	.A1N(n167),
	.A0N(\mem[8][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U280 (
	.Y(n258),
	.B1(n167),
	.B0(n366),
	.A1N(n167),
	.A0N(\mem[8][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U281 (
	.Y(n259),
	.B1(n169),
	.B0(n359),
	.A1N(n169),
	.A0N(\mem[9][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U282 (
	.Y(n260),
	.B1(n169),
	.B0(n360),
	.A1N(n169),
	.A0N(\mem[9][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U283 (
	.Y(n261),
	.B1(n169),
	.B0(n361),
	.A1N(n169),
	.A0N(\mem[9][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U284 (
	.Y(n262),
	.B1(n169),
	.B0(n362),
	.A1N(n169),
	.A0N(\mem[9][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U285 (
	.Y(n263),
	.B1(n169),
	.B0(n363),
	.A1N(n169),
	.A0N(\mem[9][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U286 (
	.Y(n264),
	.B1(n169),
	.B0(n364),
	.A1N(n169),
	.A0N(\mem[9][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U287 (
	.Y(n265),
	.B1(n169),
	.B0(n365),
	.A1N(n169),
	.A0N(\mem[9][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U288 (
	.Y(n266),
	.B1(n169),
	.B0(n366),
	.A1N(n169),
	.A0N(\mem[9][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U289 (
	.Y(n267),
	.B1(n171),
	.B0(n359),
	.A1N(n171),
	.A0N(\mem[10][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U290 (
	.Y(n268),
	.B1(n171),
	.B0(n360),
	.A1N(n171),
	.A0N(\mem[10][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U291 (
	.Y(n269),
	.B1(n171),
	.B0(n361),
	.A1N(n171),
	.A0N(\mem[10][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U292 (
	.Y(n270),
	.B1(n171),
	.B0(n362),
	.A1N(n171),
	.A0N(\mem[10][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U293 (
	.Y(n271),
	.B1(n171),
	.B0(n363),
	.A1N(n171),
	.A0N(\mem[10][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U294 (
	.Y(n272),
	.B1(n171),
	.B0(n364),
	.A1N(n171),
	.A0N(\mem[10][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U295 (
	.Y(n273),
	.B1(n171),
	.B0(n365),
	.A1N(n171),
	.A0N(\mem[10][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U296 (
	.Y(n274),
	.B1(n171),
	.B0(n366),
	.A1N(n171),
	.A0N(\mem[10][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U297 (
	.Y(n275),
	.B1(n172),
	.B0(n359),
	.A1N(n172),
	.A0N(\mem[11][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U298 (
	.Y(n276),
	.B1(n172),
	.B0(n360),
	.A1N(n172),
	.A0N(\mem[11][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U299 (
	.Y(n277),
	.B1(n172),
	.B0(n361),
	.A1N(n172),
	.A0N(\mem[11][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U300 (
	.Y(n278),
	.B1(n172),
	.B0(n362),
	.A1N(n172),
	.A0N(\mem[11][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U301 (
	.Y(n279),
	.B1(n172),
	.B0(n363),
	.A1N(n172),
	.A0N(\mem[11][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U302 (
	.Y(n280),
	.B1(n172),
	.B0(n364),
	.A1N(n172),
	.A0N(\mem[11][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U303 (
	.Y(n281),
	.B1(n172),
	.B0(n365),
	.A1N(n172),
	.A0N(\mem[11][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U304 (
	.Y(n282),
	.B1(n172),
	.B0(n366),
	.A1N(n172),
	.A0N(\mem[11][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U305 (
	.Y(n203),
	.B1(n157),
	.B0(n359),
	.A1N(n157),
	.A0N(REG2[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U306 (
	.Y(n210),
	.B1(n157),
	.B0(n366),
	.A1N(n157),
	.A0N(REG2[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U307 (
	.Y(n216),
	.B1(n159),
	.B0(n364),
	.A1N(n159),
	.A0N(REG3[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U308 (
	.Y(n283),
	.B1(n173),
	.B0(n359),
	.A1N(n173),
	.A0N(\mem[12][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U309 (
	.Y(n284),
	.B1(n173),
	.B0(n360),
	.A1N(n173),
	.A0N(\mem[12][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U310 (
	.Y(n285),
	.B1(n173),
	.B0(n361),
	.A1N(n173),
	.A0N(\mem[12][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U311 (
	.Y(n286),
	.B1(n173),
	.B0(n362),
	.A1N(n173),
	.A0N(\mem[12][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U312 (
	.Y(n287),
	.B1(n173),
	.B0(n363),
	.A1N(n173),
	.A0N(\mem[12][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U313 (
	.Y(n288),
	.B1(n173),
	.B0(n364),
	.A1N(n173),
	.A0N(\mem[12][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U314 (
	.Y(n289),
	.B1(n173),
	.B0(n365),
	.A1N(n173),
	.A0N(\mem[12][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U315 (
	.Y(n290),
	.B1(n173),
	.B0(n366),
	.A1N(n173),
	.A0N(\mem[12][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U316 (
	.Y(n291),
	.B1(n174),
	.B0(n359),
	.A1N(n174),
	.A0N(\mem[13][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U317 (
	.Y(n292),
	.B1(n174),
	.B0(n360),
	.A1N(n174),
	.A0N(\mem[13][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U318 (
	.Y(n293),
	.B1(n174),
	.B0(n361),
	.A1N(n174),
	.A0N(\mem[13][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U319 (
	.Y(n294),
	.B1(n174),
	.B0(n362),
	.A1N(n174),
	.A0N(\mem[13][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U320 (
	.Y(n295),
	.B1(n174),
	.B0(n363),
	.A1N(n174),
	.A0N(\mem[13][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U321 (
	.Y(n296),
	.B1(n174),
	.B0(n364),
	.A1N(n174),
	.A0N(\mem[13][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U322 (
	.Y(n297),
	.B1(n174),
	.B0(n365),
	.A1N(n174),
	.A0N(\mem[13][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U323 (
	.Y(n298),
	.B1(n174),
	.B0(n366),
	.A1N(n174),
	.A0N(\mem[13][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U324 (
	.Y(n299),
	.B1(n175),
	.B0(n359),
	.A1N(n175),
	.A0N(\mem[14][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U325 (
	.Y(n300),
	.B1(n175),
	.B0(n360),
	.A1N(n175),
	.A0N(\mem[14][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U326 (
	.Y(n301),
	.B1(n175),
	.B0(n361),
	.A1N(n175),
	.A0N(\mem[14][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U327 (
	.Y(n302),
	.B1(n175),
	.B0(n362),
	.A1N(n175),
	.A0N(\mem[14][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U328 (
	.Y(n303),
	.B1(n175),
	.B0(n363),
	.A1N(n175),
	.A0N(\mem[14][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U329 (
	.Y(n304),
	.B1(n175),
	.B0(n364),
	.A1N(n175),
	.A0N(\mem[14][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U330 (
	.Y(n305),
	.B1(n175),
	.B0(n365),
	.A1N(n175),
	.A0N(\mem[14][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U331 (
	.Y(n306),
	.B1(n175),
	.B0(n366),
	.A1N(n175),
	.A0N(\mem[14][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U332 (
	.Y(n307),
	.B1(n177),
	.B0(n359),
	.A1N(n177),
	.A0N(\mem[15][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U333 (
	.Y(n308),
	.B1(n177),
	.B0(n360),
	.A1N(n177),
	.A0N(\mem[15][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U334 (
	.Y(n309),
	.B1(n177),
	.B0(n361),
	.A1N(n177),
	.A0N(\mem[15][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U335 (
	.Y(n310),
	.B1(n177),
	.B0(n362),
	.A1N(n177),
	.A0N(\mem[15][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U336 (
	.Y(n311),
	.B1(n177),
	.B0(n363),
	.A1N(n177),
	.A0N(\mem[15][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U337 (
	.Y(n312),
	.B1(n177),
	.B0(n364),
	.A1N(n177),
	.A0N(\mem[15][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U338 (
	.Y(n313),
	.B1(n177),
	.B0(n365),
	.A1N(n177),
	.A0N(\mem[15][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U339 (
	.Y(n314),
	.B1(n177),
	.B0(n366),
	.A1N(n177),
	.A0N(\mem[15][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U340 (
	.Y(n219),
	.B1(n160),
	.B0(n359),
	.A1N(n160),
	.A0N(\mem[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U341 (
	.Y(n220),
	.B1(n160),
	.B0(n360),
	.A1N(n160),
	.A0N(\mem[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U342 (
	.Y(n221),
	.B1(n160),
	.B0(n361),
	.A1N(n160),
	.A0N(\mem[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U343 (
	.Y(n222),
	.B1(n160),
	.B0(n362),
	.A1N(n160),
	.A0N(\mem[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U344 (
	.Y(n223),
	.B1(n160),
	.B0(n363),
	.A1N(n160),
	.A0N(\mem[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U345 (
	.Y(n224),
	.B1(n160),
	.B0(n364),
	.A1N(n160),
	.A0N(\mem[4][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U346 (
	.Y(n225),
	.B1(n160),
	.B0(n365),
	.A1N(n160),
	.A0N(\mem[4][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U347 (
	.Y(n226),
	.B1(n160),
	.B0(n366),
	.A1N(n160),
	.A0N(\mem[4][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U348 (
	.Y(n227),
	.B1(n162),
	.B0(n359),
	.A1N(n162),
	.A0N(\mem[5][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U349 (
	.Y(n228),
	.B1(n162),
	.B0(n360),
	.A1N(n162),
	.A0N(\mem[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U350 (
	.Y(n229),
	.B1(n162),
	.B0(n361),
	.A1N(n162),
	.A0N(\mem[5][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U351 (
	.Y(n230),
	.B1(n162),
	.B0(n362),
	.A1N(n162),
	.A0N(\mem[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U352 (
	.Y(n231),
	.B1(n162),
	.B0(n363),
	.A1N(n162),
	.A0N(\mem[5][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U353 (
	.Y(n232),
	.B1(n162),
	.B0(n364),
	.A1N(n162),
	.A0N(\mem[5][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U354 (
	.Y(n233),
	.B1(n162),
	.B0(n365),
	.A1N(n162),
	.A0N(\mem[5][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U355 (
	.Y(n234),
	.B1(n162),
	.B0(n366),
	.A1N(n162),
	.A0N(\mem[5][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U356 (
	.Y(n235),
	.B1(n163),
	.B0(n359),
	.A1N(n163),
	.A0N(\mem[6][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U357 (
	.Y(n236),
	.B1(n163),
	.B0(n360),
	.A1N(n163),
	.A0N(\mem[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U358 (
	.Y(n237),
	.B1(n163),
	.B0(n361),
	.A1N(n163),
	.A0N(\mem[6][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U359 (
	.Y(n238),
	.B1(n163),
	.B0(n362),
	.A1N(n163),
	.A0N(\mem[6][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U360 (
	.Y(n239),
	.B1(n163),
	.B0(n363),
	.A1N(n163),
	.A0N(\mem[6][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U361 (
	.Y(n240),
	.B1(n163),
	.B0(n364),
	.A1N(n163),
	.A0N(\mem[6][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U362 (
	.Y(n241),
	.B1(n163),
	.B0(n365),
	.A1N(n163),
	.A0N(\mem[6][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U363 (
	.Y(n242),
	.B1(n163),
	.B0(n366),
	.A1N(n163),
	.A0N(\mem[6][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U364 (
	.Y(n243),
	.B1(n166),
	.B0(n359),
	.A1N(n166),
	.A0N(\mem[7][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U365 (
	.Y(n244),
	.B1(n166),
	.B0(n360),
	.A1N(n166),
	.A0N(\mem[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U366 (
	.Y(n245),
	.B1(n166),
	.B0(n361),
	.A1N(n166),
	.A0N(\mem[7][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U367 (
	.Y(n246),
	.B1(n166),
	.B0(n362),
	.A1N(n166),
	.A0N(\mem[7][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U368 (
	.Y(n247),
	.B1(n166),
	.B0(n363),
	.A1N(n166),
	.A0N(\mem[7][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U369 (
	.Y(n248),
	.B1(n166),
	.B0(n364),
	.A1N(n166),
	.A0N(\mem[7][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U370 (
	.Y(n249),
	.B1(n166),
	.B0(n365),
	.A1N(n166),
	.A0N(\mem[7][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U371 (
	.Y(n250),
	.B1(n166),
	.B0(n366),
	.A1N(n166),
	.A0N(\mem[7][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U372 (
	.Y(n194),
	.B1(n366),
	.B0(n152),
	.A1N(n152),
	.A0N(REG0[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U373 (
	.Y(n202),
	.B1(n155),
	.B0(n366),
	.A1N(n155),
	.A0N(REG1[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U374 (
	.Y(n195),
	.B1(n155),
	.B0(n359),
	.A1N(n155),
	.A0N(REG1[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U375 (
	.Y(n358),
	.A(WrEn), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U376 (
	.Y(n178),
	.B0(n357),
	.A1(n150),
	.A0(RdData_Valid), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X4M U377 (
	.Y(n370),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X4M U378 (
	.Y(n371),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X4M U379 (
	.Y(n372),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X4M U380 (
	.Y(n373),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_test_1 (
	A, 
	B, 
	ALU_FUN, 
	Enable, 
	CLK, 
	RST, 
	ALU_OUT, 
	OUT_VALID, 
	test_si, 
	test_se, 
	gated_clk__L3_N1, 
	VDD, 
	VSS);
   input [7:0] A;
   input [7:0] B;
   input [3:0] ALU_FUN;
   input Enable;
   input CLK;
   input RST;
   output [15:0] ALU_OUT;
   output OUT_VALID;
   input test_si;
   input test_se;
   input gated_clk__L3_N1;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_OFN11_B__1_;
   wire FE_OFN7_B__5_;
   wire FE_OFN6_B__0_;
   wire N90;
   wire N91;
   wire N92;
   wire N93;
   wire N94;
   wire N95;
   wire N96;
   wire N97;
   wire N98;
   wire N99;
   wire N100;
   wire N101;
   wire N102;
   wire N103;
   wire N104;
   wire N105;
   wire N106;
   wire N107;
   wire N108;
   wire N109;
   wire N110;
   wire N111;
   wire N112;
   wire N113;
   wire N114;
   wire N115;
   wire N116;
   wire N117;
   wire N118;
   wire N119;
   wire N120;
   wire N121;
   wire N122;
   wire N123;
   wire N124;
   wire N125;
   wire N126;
   wire N127;
   wire N128;
   wire N129;
   wire N130;
   wire N131;
   wire N156;
   wire N158;
   wire n79;
   wire n83;
   wire n84;
   wire n85;
   wire n100;
   wire n101;
   wire n102;
   wire n109;
   wire n116;
   wire n123;
   wire n130;
   wire n137;
   wire n147;
   wire n150;
   wire n151;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n162;
   wire n163;
   wire n164;
   wire n165;
   wire n166;
   wire n167;
   wire n168;
   wire n169;
   wire n170;
   wire n6;
   wire n7;
   wire n8;
   wire n43;
   wire n46;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n81;
   wire n82;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n103;
   wire n104;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n148;
   wire n149;
   wire n152;
   wire n161;
   wire n171;
   wire n172;
   wire n173;
   wire n174;
   wire n175;
   wire n176;
   wire n177;
   wire n178;
   wire n179;
   wire n180;
   wire n181;
   wire n182;
   wire n183;
   wire n184;
   wire n185;
   wire n186;
   wire n187;
   wire n188;
   wire n189;
   wire n190;
   wire n191;
   wire n192;
   wire n193;
   wire n194;
   wire n195;
   wire n196;
   wire n197;
   wire n198;
   wire n199;
   wire n200;
   wire n201;
   wire n202;
   wire n203;
   wire n204;
   wire n205;
   wire n206;
   wire n207;
   wire n208;
   wire n209;
   wire n210;
   wire n211;
   wire n212;
   wire n213;
   wire n214;
   wire n215;
   wire n216;
   wire n217;
   wire n218;
   wire n219;
   wire n220;
   wire n221;
   wire n222;
   wire n223;
   wire n224;
   wire n225;
   wire n226;
   wire n227;
   wire n228;
   wire n229;
   wire n230;
   wire n231;
   wire n232;
   wire n233;
   wire n234;
   wire n235;
   wire n236;
   wire n237;
   wire n238;
   wire n239;
   wire n240;
   wire n241;
   wire n242;
   wire n243;
   wire n244;
   wire n245;
   wire n246;
   wire n247;
   wire n248;
   wire n249;
   wire n250;
   wire n251;
   wire n252;
   wire n253;
   wire n254;
   wire n258;
   wire n259;
   wire [7:0] A_;
   wire [7:0] B_;

   // Module instantiations
   BUFX4M FE_OFC11_B__1_ (
	.Y(FE_OFN11_B__1_),
	.A(B_[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX6M FE_OFC7_B__5_ (
	.Y(FE_OFN7_B__5_),
	.A(B_[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX10M FE_OFC6_B__0_ (
	.Y(FE_OFN6_B__0_),
	.A(B_[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX4M \B__reg[7]  (
	.SI(B_[6]),
	.SE(test_se),
	.RN(RST),
	.Q(B_[7]),
	.D(B[7]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M OUT_VALID_reg (
	.SI(n177),
	.SE(test_se),
	.RN(RST),
	.Q(OUT_VALID),
	.D(Enable),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[7]  (
	.SI(ALU_OUT[6]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[7]),
	.D(n169),
	.CK(gated_clk__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[6]  (
	.SI(ALU_OUT[5]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[6]),
	.D(n168),
	.CK(gated_clk__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[5]  (
	.SI(ALU_OUT[4]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[5]),
	.D(n167),
	.CK(gated_clk__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[3]  (
	.SI(ALU_OUT[2]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[3]),
	.D(n165),
	.CK(gated_clk__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[2]  (
	.SI(ALU_OUT[1]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[2]),
	.D(n164),
	.CK(gated_clk__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[8]  (
	.SI(ALU_OUT[7]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[8]),
	.D(n170),
	.CK(gated_clk__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[15]  (
	.SI(ALU_OUT[14]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[15]),
	.D(n246),
	.CK(gated_clk__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[14]  (
	.SI(ALU_OUT[13]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[14]),
	.D(n247),
	.CK(gated_clk__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[13]  (
	.SI(ALU_OUT[12]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[13]),
	.D(n248),
	.CK(gated_clk__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[12]  (
	.SI(ALU_OUT[11]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[12]),
	.D(n249),
	.CK(gated_clk__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[11]  (
	.SI(ALU_OUT[10]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[11]),
	.D(n250),
	.CK(gated_clk__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[10]  (
	.SI(ALU_OUT[9]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[10]),
	.D(n251),
	.CK(gated_clk__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[9]  (
	.SI(ALU_OUT[8]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[9]),
	.D(n252),
	.CK(gated_clk__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \A__reg[2]  (
	.SI(n93),
	.SE(test_se),
	.RN(RST),
	.Q(A_[2]),
	.D(A[2]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \A__reg[1]  (
	.SI(n92),
	.SE(test_se),
	.RN(RST),
	.Q(A_[1]),
	.D(A[1]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \A__reg[0]  (
	.SI(ALU_OUT[15]),
	.SE(test_se),
	.RN(RST),
	.Q(A_[0]),
	.D(A[0]),
	.CK(gated_clk__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \A__reg[3]  (
	.SI(n229),
	.SE(test_se),
	.RN(RST),
	.Q(A_[3]),
	.D(A[3]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX1M \A__reg[4]  (
	.SI(n209),
	.SE(n259),
	.RN(RST),
	.Q(A_[4]),
	.D(A[4]),
	.CK(gated_clk__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX2M \B__reg[6]  (
	.SI(FE_OFN7_B__5_),
	.SE(test_se),
	.RN(RST),
	.Q(B_[6]),
	.D(B[6]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \A__reg[6]  (
	.SI(A_[5]),
	.SE(test_se),
	.RN(RST),
	.Q(A_[6]),
	.D(A[6]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX1M \ALU_OUT_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[0]),
	.D(n162),
	.CK(gated_clk__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX1M \ALU_OUT_reg[4]  (
	.SI(ALU_OUT[3]),
	.SE(n259),
	.RN(RST),
	.Q(ALU_OUT[4]),
	.D(n166),
	.CK(gated_clk__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX1M \ALU_OUT_reg[1]  (
	.SI(ALU_OUT[0]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[1]),
	.D(n163),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX1M \B__reg[3]  (
	.SI(n228),
	.SE(test_se),
	.RN(RST),
	.Q(B_[3]),
	.D(B[3]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \B__reg[1]  (
	.SI(n94),
	.SE(test_se),
	.RN(RST),
	.Q(B_[1]),
	.D(B[1]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX2M \B__reg[4]  (
	.SI(n211),
	.SE(test_se),
	.RN(RST),
	.Q(B_[4]),
	.D(B[4]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX1M \B__reg[2]  (
	.SI(FE_OFN11_B__1_),
	.SE(test_se),
	.RN(RST),
	.Q(B_[2]),
	.D(B[2]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \A__reg[5]  (
	.SI(n200),
	.SE(test_se),
	.RN(RST),
	.Q(A_[5]),
	.D(A[5]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX2M \B__reg[5]  (
	.SI(n199),
	.SE(test_se),
	.RN(RST),
	.Q(B_[5]),
	.D(B[5]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX2M \B__reg[0]  (
	.SI(n176),
	.SE(test_se),
	.RN(RST),
	.Q(B_[0]),
	.D(B[0]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX8M \A__reg[7]  (
	.SI(n183),
	.SE(test_se),
	.RN(RST),
	.Q(A_[7]),
	.D(A[7]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U49 (
	.Y(n6),
	.A(B_[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U50 (
	.Y(n7),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U51 (
	.Y(n8),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U53 (
	.Y(n43),
	.B(Enable),
	.A(n225), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U56 (
	.Y(n46),
	.B(n43),
	.A(N124), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U57 (
	.Y(n162),
	.B(n135),
	.A(n46), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX1M U58 (
	.Y(n136),
	.C(n118),
	.B(n53),
	.AN(n244), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U59 (
	.Y(n135),
	.B1(Enable),
	.B0(ALU_OUT[0]),
	.A1N(n134),
	.A0(n133), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BXLM U61 (
	.Y(n88),
	.B(A_[5]),
	.AN(FE_OFN7_B__5_), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2BB1XLM U62 (
	.Y(n81),
	.B0(FE_OFN11_B__1_),
	.A1N(n82),
	.A0N(A_[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR2XLM U64 (
	.Y(n55),
	.B(A_[6]),
	.A(B_[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BXLM U65 (
	.Y(n184),
	.B(B_[6]),
	.AN(n183), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U66 (
	.Y(n163),
	.S0(Enable),
	.B(n171),
	.A(ALU_OUT[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211XLM U68 (
	.Y(n198),
	.C0(n193),
	.B0(n194),
	.A1(n224),
	.A0(A_[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U69 (
	.Y(n225),
	.A(n136), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U70 (
	.Y(n232),
	.A(n213), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U71 (
	.Y(n146),
	.A(n85), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U72 (
	.Y(n253),
	.A(n150), 
	.VDD(VDD), 
	.VSS(VSS));
   OA21X2M U73 (
	.Y(n174),
	.B0(n79),
	.A1(n172),
	.A0(n173), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U74 (
	.Y(n213),
	.B0(n54),
	.A1(n242),
	.A0(n124), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U75 (
	.Y(n226),
	.A(n112), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX2M U76 (
	.Y(n112),
	.C(n242),
	.B(n147),
	.AN(n244), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U77 (
	.Y(n241),
	.A(n121), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U78 (
	.Y(n214),
	.A(n231), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U79 (
	.Y(n208),
	.A(n233), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U80 (
	.Y(n223),
	.A(n138), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U81 (
	.Y(n230),
	.A(n212), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U82 (
	.Y(n124),
	.A(n101), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U84 (
	.Y(n178),
	.B1(n241),
	.B0(N115),
	.A1(n226),
	.A0(N106), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U85 (
	.Y(n186),
	.C(n51),
	.B(n50),
	.A(n49), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U86 (
	.Y(n49),
	.S0(n184),
	.B(n230),
	.A(n231), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U87 (
	.Y(n50),
	.S0(n185),
	.B(n232),
	.A(n233), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U88 (
	.Y(n51),
	.B1(n241),
	.B0(N114),
	.A1(n55),
	.A0(n79), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4BX1M U89 (
	.Y(n85),
	.D(ALU_FUN[0]),
	.C(n101),
	.B(n242),
	.AN(N158), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U90 (
	.Y(n235),
	.B1(n241),
	.B0(N110),
	.A1(n234),
	.A0(n79), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U91 (
	.Y(n150),
	.B(Enable),
	.A(n113), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U92 (
	.Y(n113),
	.B0(n212),
	.A1(n226),
	.A0(N107), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U93 (
	.Y(n128),
	.A(n83), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U94 (
	.Y(n83),
	.B0(n85),
	.A2(n84),
	.A1(ALU_FUN[1]),
	.A0(N156), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U95 (
	.Y(n84),
	.C(ALU_FUN[0]),
	.B(ALU_FUN[2]),
	.A(n242), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X2M U96 (
	.Y(n143),
	.C(n245),
	.B(ALU_FUN[0]),
	.A(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U97 (
	.Y(n100),
	.C(n242),
	.B(ALU_FUN[2]),
	.A(n243), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U98 (
	.Y(n196),
	.B1(n227),
	.B0(N95),
	.A1(n226),
	.A0(N104), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U99 (
	.Y(n145),
	.C1(n226),
	.C0(N100),
	.B1(n227),
	.B0(N91),
	.A1(n241),
	.A0(N109), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U100 (
	.Y(n172),
	.A(n110), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U101 (
	.Y(n173),
	.A(n108), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U102 (
	.Y(n180),
	.S0(n52),
	.B(n231),
	.A(n230), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U103 (
	.Y(n52),
	.B(n176),
	.A(n177), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX2M U104 (
	.Y(n233),
	.C(n53),
	.B(ALU_FUN[2]),
	.AN(ALU_FUN[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX2M U105 (
	.Y(n231),
	.C(n124),
	.B(ALU_FUN[0]),
	.AN(ALU_FUN[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U106 (
	.Y(n147),
	.B(ALU_FUN[1]),
	.A(ALU_FUN[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX2M U107 (
	.Y(n138),
	.C(n124),
	.B(ALU_FUN[0]),
	.AN(n242), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U108 (
	.Y(n212),
	.B0(n54),
	.A1(ALU_FUN[2]),
	.A0(n53), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX2M U109 (
	.Y(n121),
	.C(n118),
	.B(n53),
	.AN(ALU_FUN[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U110 (
	.Y(n242),
	.A(ALU_FUN[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X2M U111 (
	.Y(n79),
	.C(n244),
	.B(ALU_FUN[3]),
	.A(n147), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U112 (
	.Y(n227),
	.A(n115), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX2M U113 (
	.Y(n115),
	.C(n244),
	.B(n147),
	.AN(ALU_FUN[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U114 (
	.Y(n101),
	.B(n118),
	.A(ALU_FUN[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U115 (
	.Y(n254),
	.A(Enable), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U116 (
	.Y(n154),
	.B(Enable),
	.A(n241), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U117 (
	.Y(n224),
	.A(n114), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BX1M U118 (
	.Y(n114),
	.D(ALU_FUN[3]),
	.C(ALU_FUN[2]),
	.B(ALU_FUN[1]),
	.AN(ALU_FUN[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U119 (
	.Y(n244),
	.A(ALU_FUN[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U120 (
	.Y(n118),
	.A(ALU_FUN[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U122 (
	.Y(n243),
	.A(ALU_FUN[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U123 (
	.Y(n53),
	.B(n243),
	.A(ALU_FUN[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X2M U124 (
	.Y(n54),
	.C(n147),
	.B(ALU_FUN[3]),
	.A(ALU_FUN[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22XLM U125 (
	.Y(n161),
	.B1(n223),
	.B0(A_[2]),
	.A1(n225),
	.A0(N125), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U126 (
	.Y(n92),
	.A(A_[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U127 (
	.Y(n93),
	.A(A_[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X2M U128 (
	.Y(n103),
	.C0(n60),
	.B0(n56),
	.A1(n98),
	.A0(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U129 (
	.Y(n99),
	.B0(n61),
	.A2(n95),
	.A1(n96),
	.A0(n97), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U130 (
	.Y(n95),
	.B0(A_[1]),
	.A1(n94),
	.A0(A_[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U131 (
	.Y(n97),
	.A(n234), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI31X1M U132 (
	.Y(n87),
	.B0(n98),
	.A2(n56),
	.A1(n57),
	.A0(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X2M U133 (
	.Y(n86),
	.C0(n234),
	.B0(n81),
	.A1(n82),
	.A0(A_[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U134 (
	.Y(N158),
	.B0(n172),
	.A1(n108),
	.A0(n91), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X2M U135 (
	.Y(n90),
	.C0(n104),
	.B0(n55),
	.A1(n105),
	.A0(n89), 
	.VDD(VDD), 
	.VSS(VSS));
   OA22X2M U136 (
	.Y(n89),
	.B1(n199),
	.B0(A_[4]),
	.A1(n87),
	.A0(n60), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U137 (
	.Y(n133),
	.C(n129),
	.B(n131),
	.A(n132), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U138 (
	.Y(n132),
	.S0(A_[0]),
	.B(n126),
	.A(n127), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U139 (
	.Y(n129),
	.B(n227),
	.A(N90), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U140 (
	.Y(n131),
	.B0(n128),
	.A1(n226),
	.A0(N99), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U141 (
	.Y(n202),
	.B1(n241),
	.B0(N112),
	.A1(n60),
	.A0(n79), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U142 (
	.Y(n234),
	.B(n61),
	.A(n57), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U143 (
	.Y(n218),
	.B1(n227),
	.B0(N93),
	.A1(n226),
	.A0(N102), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U144 (
	.Y(n245),
	.B0(n173),
	.A1(n110),
	.A0(n111), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U145 (
	.Y(n106),
	.A(n105), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X2M U146 (
	.Y(n107),
	.C0(n103),
	.B0(n104),
	.A1(n199),
	.A0(A_[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U147 (
	.Y(n219),
	.B0(n217),
	.A1(n241),
	.A0(N111), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U148 (
	.Y(n217),
	.S0(A_[3]),
	.B(n215),
	.A(n216), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U149 (
	.Y(n216),
	.B(n211),
	.A(n212), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U150 (
	.Y(n82),
	.B(n94),
	.A(A_[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U151 (
	.Y(n56),
	.B(n211),
	.A(A_[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U152 (
	.Y(n229),
	.A(A_[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U153 (
	.Y(n57),
	.B(n228),
	.A(A_[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U154 (
	.Y(n179),
	.S0(n58),
	.B(n233),
	.A(n232), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2XLM U155 (
	.Y(n58),
	.B(A_[7]),
	.A(B_[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U156 (
	.Y(n108),
	.B(n176),
	.A(B_[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U157 (
	.Y(n105),
	.B(FE_OFN7_B__5_),
	.AN(A_[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U158 (
	.Y(n140),
	.S0(FE_OFN11_B__1_),
	.B(n213),
	.A(n79), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X1M U159 (
	.Y(n190),
	.S0(FE_OFN7_B__5_),
	.B(n213),
	.A(n79), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U160 (
	.Y(n144),
	.S0(A_[1]),
	.B(n141),
	.A(n142), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U161 (
	.Y(n142),
	.B(n139),
	.A(n208), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U162 (
	.Y(n141),
	.B(n140),
	.A(n214), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U163 (
	.Y(n139),
	.S0(FE_OFN11_B__1_),
	.B(n79),
	.A(n212), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U164 (
	.Y(n177),
	.A(B_[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U165 (
	.Y(n193),
	.S0(A_[5]),
	.B(n191),
	.A(n192), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U166 (
	.Y(n192),
	.B(n189),
	.A(n208), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U167 (
	.Y(n191),
	.B(n190),
	.A(n214), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X1M U168 (
	.Y(n189),
	.S0(FE_OFN7_B__5_),
	.B(n79),
	.A(n212), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U169 (
	.Y(n209),
	.A(A_[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U170 (
	.Y(n104),
	.A(n88), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U171 (
	.Y(n183),
	.A(A_[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B11X2M U172 (
	.Y(n120),
	.C0(n119),
	.B0(Enable),
	.A1N(A_[1]),
	.A0(n138), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U173 (
	.Y(n127),
	.B(n122),
	.AN(n208), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U174 (
	.Y(n126),
	.B(n125),
	.AN(n214), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X1M U175 (
	.Y(n195),
	.S0(FE_OFN7_B__5_),
	.B(n214),
	.A(n208), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U176 (
	.Y(n148),
	.S0(FE_OFN11_B__1_),
	.B(n231),
	.A(n233), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U177 (
	.Y(n204),
	.S0(n201),
	.B(n230),
	.A(n231), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U178 (
	.Y(n201),
	.B(n199),
	.A(n200), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U179 (
	.Y(n200),
	.A(A_[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OA21X2M U180 (
	.Y(n210),
	.B0(n208),
	.A1(n211),
	.A0(n209), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U181 (
	.Y(n237),
	.S0(n59),
	.B(n231),
	.A(n230), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U182 (
	.Y(n59),
	.B(n228),
	.A(n229), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2B1X1M U184 (
	.Y(n134),
	.B0(n120),
	.A1N(n121),
	.A0(N108), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX2M U185 (
	.Y(n171),
	.C(n149),
	.B(n152),
	.AN(n161), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X2M U186 (
	.Y(n152),
	.C0(n143),
	.B0(n144),
	.A1(n224),
	.A0(A_[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X2M U187 (
	.Y(n149),
	.C(n145),
	.B(n146),
	.A(n148), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U189 (
	.Y(n164),
	.B0(n102),
	.A1(n254),
	.A0(ALU_OUT[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U190 (
	.Y(n102),
	.B0(n254),
	.A2(n238),
	.A1(n239),
	.A0(n240), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U191 (
	.Y(n239),
	.B1(n226),
	.B0(N101),
	.A1(n227),
	.A0(N92), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X2M U192 (
	.Y(n238),
	.C(n235),
	.B(n236),
	.A(n237), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U195 (
	.Y(n248),
	.A(n158), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U196 (
	.Y(n158),
	.C0(n253),
	.B1(n154),
	.B0(N121),
	.A1(n254),
	.A0(ALU_OUT[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U197 (
	.Y(n247),
	.A(n159), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U198 (
	.Y(n159),
	.C0(n253),
	.B1(n154),
	.B0(N122),
	.A1(n254),
	.A0(ALU_OUT[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U199 (
	.Y(n246),
	.A(n160), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U200 (
	.Y(n160),
	.C0(n253),
	.B1(n154),
	.B0(N123),
	.A1(n254),
	.A0(ALU_OUT[15]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22XLM U201 (
	.Y(n221),
	.B1(n8),
	.B0(n214),
	.A1(n225),
	.A0(N127), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U202 (
	.Y(n252),
	.A(n153), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U203 (
	.Y(n153),
	.C0(n253),
	.B1(n154),
	.B0(N117),
	.A1(n254),
	.A0(ALU_OUT[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U204 (
	.Y(n165),
	.B0(n109),
	.A1(n254),
	.A0(ALU_OUT[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U205 (
	.Y(n109),
	.B0(n254),
	.A2(n220),
	.A1(n221),
	.A0(n222), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U206 (
	.Y(n222),
	.C0(n210),
	.B1(n224),
	.B0(A_[2]),
	.A1(n223),
	.A0(A_[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X2M U207 (
	.Y(n220),
	.C0(n218),
	.B0(n219),
	.A1(n79),
	.A0(n56), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B11X2M U208 (
	.Y(n170),
	.C0(n150),
	.B0(n151),
	.A1N(Enable),
	.A0(n117), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U209 (
	.Y(n151),
	.B(n254),
	.A(ALU_OUT[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U210 (
	.Y(n251),
	.A(n155), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U211 (
	.Y(n155),
	.C0(n253),
	.B1(n154),
	.B0(N118),
	.A1(n254),
	.A0(ALU_OUT[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U212 (
	.Y(n250),
	.A(n156), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U213 (
	.Y(n156),
	.C0(n253),
	.B1(n154),
	.B0(N119),
	.A1(n254),
	.A0(ALU_OUT[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U214 (
	.Y(n249),
	.A(n157), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U215 (
	.Y(n157),
	.C0(n253),
	.B1(n154),
	.B0(N120),
	.A1(n254),
	.A0(ALU_OUT[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U216 (
	.Y(n166),
	.B0(n116),
	.A1(n254),
	.A0(ALU_OUT[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U217 (
	.Y(n116),
	.B0(n254),
	.A2(n205),
	.A1(n206),
	.A0(n207), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U218 (
	.Y(n206),
	.B1(n226),
	.B0(N103),
	.A1(n227),
	.A0(N94), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X2M U219 (
	.Y(n205),
	.C(n202),
	.B(n203),
	.A(n204), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U220 (
	.Y(n169),
	.B0(n137),
	.A1(n254),
	.A0(ALU_OUT[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U221 (
	.Y(n137),
	.B0(n254),
	.A1(n181),
	.A0(n182), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X2M U222 (
	.Y(n181),
	.C(n178),
	.B(n179),
	.A(n180), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U223 (
	.Y(n168),
	.B0(n130),
	.A1(n254),
	.A0(ALU_OUT[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U224 (
	.Y(n130),
	.B0(n254),
	.A2(n186),
	.A1(n187),
	.A0(n188), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U225 (
	.Y(n187),
	.B1(n226),
	.B0(N105),
	.A1(n227),
	.A0(N96), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U226 (
	.Y(n167),
	.B0(n123),
	.A1(n254),
	.A0(ALU_OUT[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U227 (
	.Y(n123),
	.B0(n254),
	.A1(n197),
	.A0(n198), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X2M U228 (
	.Y(n197),
	.C0(n195),
	.B0(n196),
	.A1(n241),
	.A0(N113), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U229 (
	.Y(n211),
	.A(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U230 (
	.Y(n228),
	.A(B_[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR2XLM U231 (
	.Y(n60),
	.B(A_[4]),
	.A(B_[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2XLM U232 (
	.Y(n61),
	.B(n229),
	.A(B_[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U233 (
	.Y(n199),
	.A(B_[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U234 (
	.Y(n98),
	.B(n209),
	.A(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U235 (
	.Y(n215),
	.B(n62),
	.AN(n214), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2XLM U236 (
	.Y(n62),
	.S0(n8),
	.B(n213),
	.A(n79), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U237 (
	.Y(n236),
	.S0(n63),
	.B(n233),
	.A(n232), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2XLM U238 (
	.Y(n63),
	.B(B_[2]),
	.A(A_[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U239 (
	.Y(n203),
	.S0(n64),
	.B(n233),
	.A(n232), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2XLM U240 (
	.Y(n64),
	.B(A_[4]),
	.A(B_[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U241 (
	.Y(n185),
	.B(A_[6]),
	.A(B_[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI32XLM U242 (
	.Y(n111),
	.B1(n183),
	.B0(B_[6]),
	.A2(n55),
	.A1(n106),
	.A0(n107), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U243 (
	.Y(n91),
	.B0(n90),
	.A1(n183),
	.A0(B_[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U244 (
	.Y(n110),
	.B(n177),
	.A(A_[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U245 (
	.Y(n176),
	.A(A_[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2XLM U246 (
	.Y(n119),
	.S0(FE_OFN6_B__0_),
	.B(n214),
	.A(n208), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2XLM U247 (
	.Y(n122),
	.S0(FE_OFN6_B__0_),
	.B(n79),
	.A(n212), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2XLM U248 (
	.Y(n125),
	.S0(FE_OFN6_B__0_),
	.B(n213),
	.A(n79), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U249 (
	.Y(n94),
	.A(FE_OFN6_B__0_), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U250 (
	.Y(n194),
	.B1(n223),
	.B0(A_[6]),
	.A1(n225),
	.A0(N129), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222XLM U251 (
	.Y(n240),
	.C1(n223),
	.C0(A_[3]),
	.B1(n224),
	.B0(A_[1]),
	.A1(n225),
	.A0(N126), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X2M U252 (
	.Y(n182),
	.C0(n174),
	.B0(n175),
	.A1(n224),
	.A0(A_[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI31XLM U253 (
	.Y(n96),
	.B0(FE_OFN11_B__1_),
	.A2(n92),
	.A1(n93),
	.A0(FE_OFN6_B__0_), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22XLM U254 (
	.Y(n175),
	.B1(n225),
	.B0(N131),
	.A1(n227),
	.A0(N97), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222XLM U255 (
	.Y(n117),
	.C1(n227),
	.C0(N98),
	.B1(n224),
	.B0(A_[7]),
	.A1(n241),
	.A0(N116), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222XLM U256 (
	.Y(n188),
	.C1(n223),
	.C0(A_[7]),
	.B1(n224),
	.B0(A_[5]),
	.A1(n225),
	.A0(N130), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U257 (
	.Y(n207),
	.C1(n223),
	.C0(A_[5]),
	.B1(n224),
	.B0(A_[3]),
	.A1(n225),
	.A0(N128), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U258 (
	.Y(N156),
	.B(n245),
	.A(N158), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U260 (
	.Y(n258),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U261 (
	.Y(n259),
	.A(n258), 
	.VDD(VDD), 
	.VSS(VSS));
   ALU_DW01_sub_0 sub_34 (
	.A({ 1'b0,
		A_[7],
		A_[6],
		A_[5],
		A_[4],
		A_[3],
		A_[2],
		A_[1],
		A_[0] }),
	.B({ 1'b0,
		B_[7],
		B_[6],
		FE_OFN7_B__5_,
		B_[4],
		n8,
		B_[2],
		FE_OFN11_B__1_,
		FE_OFN6_B__0_ }),
	.CI(1'b0),
	.DIFF({ N107,
		N106,
		N105,
		N104,
		N103,
		N102,
		N101,
		N100,
		N99 }),
	.n94(n94),
	.n228(n228),
	.n199(n199),
	.n211(n211),
	.n92(n92),
	.n177(n177), 
	.VDD(VDD), 
	.VSS(VSS));
   ALU_DW01_add_0 add_33 (
	.A({ 1'b0,
		A_[7],
		A_[6],
		A_[5],
		A_[4],
		A_[3],
		A_[2],
		A_[1],
		A_[0] }),
	.B({ 1'b0,
		B_[7],
		B_[6],
		FE_OFN7_B__5_,
		B_[4],
		n8,
		B_[2],
		FE_OFN11_B__1_,
		FE_OFN6_B__0_ }),
	.CI(1'b0),
	.SUM({ N98,
		N97,
		N96,
		N95,
		N94,
		N93,
		N92,
		N91,
		N90 }),
	.n92(n92), 
	.VDD(VDD), 
	.VSS(VSS));
   ALU_DW02_mult_0 mult_35 (
	.A({ A_[7],
		A_[6],
		A_[5],
		A_[4],
		A_[3],
		A_[2],
		A_[1],
		A_[0] }),
	.B({ B_[7],
		B_[6],
		FE_OFN7_B__5_,
		B_[4],
		n8,
		B_[2],
		FE_OFN11_B__1_,
		FE_OFN6_B__0_ }),
	.TC(1'b0),
	.PRODUCT({ N123,
		N122,
		N121,
		N120,
		N119,
		N118,
		N117,
		N116,
		N115,
		N114,
		N113,
		N112,
		N111,
		N110,
		N109,
		N108 }),
	.n200(n200),
	.n183(n183),
	.n209(n209),
	.n92(n92),
	.n93(n93),
	.n229(n229),
	.n177(n177), 
	.VDD(VDD), 
	.VSS(VSS));
   ALU_DW_div_uns_1 div_36 (
	.a({ A_[7],
		A_[6],
		A_[5],
		A_[4],
		A_[3],
		A_[2],
		A_[1],
		A_[0] }),
	.b({ B_[7],
		B_[6],
		FE_OFN7_B__5_,
		B_[4],
		n7,
		B_[2],
		FE_OFN11_B__1_,
		FE_OFN6_B__0_ }),
	.quotient({ N131,
		N130,
		N129,
		N128,
		N127,
		N126,
		N125,
		N124 }),
	.n200(n200),
	.n209(n209),
	.FE_PT1_n92(n92),
	.FE_PT1_n93(n93),
	.n176(n176),
	.n183(n183),
	.n177(n177), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_DW01_sub_0 (
	A, 
	B, 
	CI, 
	DIFF, 
	CO, 
	n94, 
	n228, 
	n199, 
	n211, 
	n92, 
	n177, 
	VDD, 
	VSS);
   input [8:0] A;
   input [8:0] B;
   input CI;
   output [8:0] DIFF;
   output CO;
   input n94;
   input n228;
   input n199;
   input n211;
   input n92;
   input n177;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n3;
   wire n4;
   wire n8;
   wire [9:0] carry;

   // Module instantiations
   ADDFX2M U2_4 (
	.S(DIFF[4]),
	.CO(carry[5]),
	.CI(carry[4]),
	.B(n199),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_2 (
	.S(DIFF[2]),
	.CO(carry[3]),
	.CI(carry[2]),
	.B(n228),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_3 (
	.S(DIFF[3]),
	.CO(carry[4]),
	.CI(carry[3]),
	.B(n211),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_6 (
	.S(DIFF[6]),
	.CO(carry[7]),
	.CI(carry[6]),
	.B(n3),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_1 (
	.S(DIFF[1]),
	.CO(carry[2]),
	.CI(carry[1]),
	.B(n8),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_5 (
	.S(DIFF[5]),
	.CO(carry[6]),
	.CI(carry[5]),
	.B(n4),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_7 (
	.S(DIFF[7]),
	.CO(carry[8]),
	.CI(carry[7]),
	.B(n177),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U2 (
	.Y(n4),
	.A(B[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U3 (
	.Y(n8),
	.A(B[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U4 (
	.Y(carry[1]),
	.B(n92),
	.A(B[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U6 (
	.Y(DIFF[0]),
	.B(A[0]),
	.A(n94), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U10 (
	.Y(n3),
	.A(B[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U12 (
	.Y(DIFF[8]),
	.A(carry[8]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_DW01_add_0 (
	A, 
	B, 
	CI, 
	SUM, 
	CO, 
	n92, 
	VDD, 
	VSS);
   input [8:0] A;
   input [8:0] B;
   input CI;
   output [8:0] SUM;
   output CO;
   input n92;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n3;
   wire [8:1] carry;

   // Module instantiations
   ADDFX2M U1_6 (
	.S(SUM[6]),
	.CO(carry[7]),
	.CI(carry[6]),
	.B(B[6]),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.CI(carry[4]),
	.B(B[4]),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.CI(carry[2]),
	.B(B[2]),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.CI(carry[3]),
	.B(B[3]),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.CI(carry[5]),
	.B(B[5]),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.CI(carry[1]),
	.B(B[1]),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_7 (
	.S(SUM[7]),
	.CO(SUM[8]),
	.CI(carry[7]),
	.B(B[7]),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U2 (
	.Y(SUM[0]),
	.B(n92),
	.A(B[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U3 (
	.Y(n3),
	.B(A[0]),
	.A(B[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U4 (
	.Y(carry[1]),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_DW02_mult_0 (
	A, 
	B, 
	TC, 
	PRODUCT, 
	n200, 
	n183, 
	n209, 
	n92, 
	n93, 
	n229, 
	n177, 
	VDD, 
	VSS);
   input [7:0] A;
   input [7:0] B;
   input TC;
   output [15:0] PRODUCT;
   input n200;
   input n183;
   input n209;
   input n92;
   input n93;
   input n229;
   input n177;
   inout VDD;
   inout VSS;

   // Internal wires
   wire \ab[7][7] ;
   wire \ab[7][6] ;
   wire \ab[7][5] ;
   wire \ab[7][4] ;
   wire \ab[7][3] ;
   wire \ab[7][2] ;
   wire \ab[7][1] ;
   wire \ab[7][0] ;
   wire \ab[6][7] ;
   wire \ab[6][6] ;
   wire \ab[6][5] ;
   wire \ab[6][4] ;
   wire \ab[6][3] ;
   wire \ab[6][2] ;
   wire \ab[6][1] ;
   wire \ab[6][0] ;
   wire \ab[5][7] ;
   wire \ab[5][6] ;
   wire \ab[5][5] ;
   wire \ab[5][4] ;
   wire \ab[5][3] ;
   wire \ab[5][2] ;
   wire \ab[5][1] ;
   wire \ab[5][0] ;
   wire \ab[4][7] ;
   wire \ab[4][6] ;
   wire \ab[4][5] ;
   wire \ab[4][4] ;
   wire \ab[4][3] ;
   wire \ab[4][2] ;
   wire \ab[4][1] ;
   wire \ab[4][0] ;
   wire \ab[3][7] ;
   wire \ab[3][6] ;
   wire \ab[3][5] ;
   wire \ab[3][4] ;
   wire \ab[3][3] ;
   wire \ab[3][2] ;
   wire \ab[3][1] ;
   wire \ab[3][0] ;
   wire \ab[2][7] ;
   wire \ab[2][6] ;
   wire \ab[2][5] ;
   wire \ab[2][4] ;
   wire \ab[2][3] ;
   wire \ab[2][2] ;
   wire \ab[2][1] ;
   wire \ab[2][0] ;
   wire \ab[1][7] ;
   wire \ab[1][6] ;
   wire \ab[1][5] ;
   wire \ab[1][4] ;
   wire \ab[1][3] ;
   wire \ab[1][2] ;
   wire \ab[1][1] ;
   wire \ab[1][0] ;
   wire \ab[0][7] ;
   wire \ab[0][6] ;
   wire \ab[0][5] ;
   wire \ab[0][4] ;
   wire \ab[0][3] ;
   wire \ab[0][2] ;
   wire \ab[0][1] ;
   wire \CARRYB[7][6] ;
   wire \CARRYB[7][5] ;
   wire \CARRYB[7][4] ;
   wire \CARRYB[7][3] ;
   wire \CARRYB[7][2] ;
   wire \CARRYB[7][1] ;
   wire \CARRYB[7][0] ;
   wire \CARRYB[6][6] ;
   wire \CARRYB[6][5] ;
   wire \CARRYB[6][4] ;
   wire \CARRYB[6][3] ;
   wire \CARRYB[6][2] ;
   wire \CARRYB[6][1] ;
   wire \CARRYB[6][0] ;
   wire \CARRYB[5][6] ;
   wire \CARRYB[5][5] ;
   wire \CARRYB[5][4] ;
   wire \CARRYB[5][3] ;
   wire \CARRYB[5][2] ;
   wire \CARRYB[5][1] ;
   wire \CARRYB[5][0] ;
   wire \CARRYB[4][6] ;
   wire \CARRYB[4][5] ;
   wire \CARRYB[4][4] ;
   wire \CARRYB[4][3] ;
   wire \CARRYB[4][2] ;
   wire \CARRYB[4][1] ;
   wire \CARRYB[4][0] ;
   wire \CARRYB[3][6] ;
   wire \CARRYB[3][5] ;
   wire \CARRYB[3][4] ;
   wire \CARRYB[3][3] ;
   wire \CARRYB[3][2] ;
   wire \CARRYB[3][1] ;
   wire \CARRYB[3][0] ;
   wire \CARRYB[2][6] ;
   wire \CARRYB[2][5] ;
   wire \CARRYB[2][4] ;
   wire \CARRYB[2][3] ;
   wire \CARRYB[2][2] ;
   wire \CARRYB[2][1] ;
   wire \CARRYB[2][0] ;
   wire \SUMB[7][6] ;
   wire \SUMB[7][5] ;
   wire \SUMB[7][4] ;
   wire \SUMB[7][3] ;
   wire \SUMB[7][2] ;
   wire \SUMB[7][1] ;
   wire \SUMB[7][0] ;
   wire \SUMB[6][6] ;
   wire \SUMB[6][5] ;
   wire \SUMB[6][4] ;
   wire \SUMB[6][3] ;
   wire \SUMB[6][2] ;
   wire \SUMB[6][1] ;
   wire \SUMB[5][6] ;
   wire \SUMB[5][5] ;
   wire \SUMB[5][4] ;
   wire \SUMB[5][3] ;
   wire \SUMB[5][2] ;
   wire \SUMB[5][1] ;
   wire \SUMB[4][6] ;
   wire \SUMB[4][5] ;
   wire \SUMB[4][4] ;
   wire \SUMB[4][3] ;
   wire \SUMB[4][2] ;
   wire \SUMB[4][1] ;
   wire \SUMB[3][6] ;
   wire \SUMB[3][5] ;
   wire \SUMB[3][4] ;
   wire \SUMB[3][3] ;
   wire \SUMB[3][2] ;
   wire \SUMB[3][1] ;
   wire \SUMB[2][6] ;
   wire \SUMB[2][5] ;
   wire \SUMB[2][4] ;
   wire \SUMB[2][3] ;
   wire \SUMB[2][2] ;
   wire \SUMB[2][1] ;
   wire \SUMB[1][6] ;
   wire \SUMB[1][5] ;
   wire \SUMB[1][4] ;
   wire \SUMB[1][3] ;
   wire \SUMB[1][2] ;
   wire \SUMB[1][1] ;
   wire \A1[12] ;
   wire \A1[11] ;
   wire \A1[10] ;
   wire \A1[9] ;
   wire \A1[8] ;
   wire \A1[7] ;
   wire \A1[6] ;
   wire \A1[4] ;
   wire \A1[3] ;
   wire \A1[2] ;
   wire \A1[1] ;
   wire \A1[0] ;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n27;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;

   // Module instantiations
   ADDFX2M S2_6_2 (
	.S(\SUMB[6][2] ),
	.CO(\CARRYB[6][2] ),
	.CI(\SUMB[5][3] ),
	.B(\CARRYB[5][2] ),
	.A(\ab[6][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_5_3 (
	.S(\SUMB[5][3] ),
	.CO(\CARRYB[5][3] ),
	.CI(\SUMB[4][4] ),
	.B(\CARRYB[4][3] ),
	.A(\ab[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_5_2 (
	.S(\SUMB[5][2] ),
	.CO(\CARRYB[5][2] ),
	.CI(\SUMB[4][3] ),
	.B(\CARRYB[4][2] ),
	.A(\ab[5][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_4_4 (
	.S(\SUMB[4][4] ),
	.CO(\CARRYB[4][4] ),
	.CI(\SUMB[3][5] ),
	.B(\CARRYB[3][4] ),
	.A(\ab[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_4_2 (
	.S(\SUMB[4][2] ),
	.CO(\CARRYB[4][2] ),
	.CI(\SUMB[3][3] ),
	.B(\CARRYB[3][2] ),
	.A(\ab[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_3_4 (
	.S(\SUMB[3][4] ),
	.CO(\CARRYB[3][4] ),
	.CI(\SUMB[2][5] ),
	.B(\CARRYB[2][4] ),
	.A(\ab[3][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_3_2 (
	.S(\SUMB[3][2] ),
	.CO(\CARRYB[3][2] ),
	.CI(\SUMB[2][3] ),
	.B(\CARRYB[2][2] ),
	.A(\ab[3][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_2_2 (
	.S(\SUMB[2][2] ),
	.CO(\CARRYB[2][2] ),
	.CI(\SUMB[1][3] ),
	.B(n6),
	.A(\ab[2][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_6_4 (
	.S(\SUMB[6][4] ),
	.CO(\CARRYB[6][4] ),
	.CI(\SUMB[5][5] ),
	.B(\CARRYB[5][4] ),
	.A(\ab[6][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_6_3 (
	.S(\SUMB[6][3] ),
	.CO(\CARRYB[6][3] ),
	.CI(\SUMB[5][4] ),
	.B(\CARRYB[5][3] ),
	.A(\ab[6][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_5_4 (
	.S(\SUMB[5][4] ),
	.CO(\CARRYB[5][4] ),
	.CI(\SUMB[4][5] ),
	.B(\CARRYB[4][4] ),
	.A(\ab[5][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_4_3 (
	.S(\SUMB[4][3] ),
	.CO(\CARRYB[4][3] ),
	.CI(\SUMB[3][4] ),
	.B(\CARRYB[3][3] ),
	.A(\ab[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_3_3 (
	.S(\SUMB[3][3] ),
	.CO(\CARRYB[3][3] ),
	.CI(\SUMB[2][4] ),
	.B(\CARRYB[2][3] ),
	.A(\ab[3][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_2_3 (
	.S(\SUMB[2][3] ),
	.CO(\CARRYB[2][3] ),
	.CI(\SUMB[1][4] ),
	.B(n5),
	.A(\ab[2][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_4 (
	.S(\SUMB[7][4] ),
	.CO(\CARRYB[7][4] ),
	.CI(\SUMB[6][5] ),
	.B(\CARRYB[6][4] ),
	.A(\ab[7][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_3 (
	.S(\SUMB[7][3] ),
	.CO(\CARRYB[7][3] ),
	.CI(\SUMB[6][4] ),
	.B(\CARRYB[6][3] ),
	.A(\ab[7][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_2 (
	.S(\SUMB[7][2] ),
	.CO(\CARRYB[7][2] ),
	.CI(\SUMB[6][3] ),
	.B(\CARRYB[6][2] ),
	.A(\ab[7][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_2_4 (
	.S(\SUMB[2][4] ),
	.CO(\CARRYB[2][4] ),
	.CI(\SUMB[1][5] ),
	.B(n8),
	.A(\ab[2][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S3_6_6 (
	.S(\SUMB[6][6] ),
	.CO(\CARRYB[6][6] ),
	.CI(\ab[5][7] ),
	.B(\CARRYB[5][6] ),
	.A(\ab[6][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S5_6 (
	.S(\SUMB[7][6] ),
	.CO(\CARRYB[7][6] ),
	.CI(\ab[6][7] ),
	.B(\CARRYB[6][6] ),
	.A(\ab[7][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S1_3_0 (
	.S(\A1[1] ),
	.CO(\CARRYB[3][0] ),
	.CI(\SUMB[2][1] ),
	.B(\CARRYB[2][0] ),
	.A(\ab[3][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S1_6_0 (
	.S(\A1[4] ),
	.CO(\CARRYB[6][0] ),
	.CI(\SUMB[5][1] ),
	.B(\CARRYB[5][0] ),
	.A(\ab[6][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_6_1 (
	.S(\SUMB[6][1] ),
	.CO(\CARRYB[6][1] ),
	.CI(\SUMB[5][2] ),
	.B(\CARRYB[5][1] ),
	.A(\ab[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S1_5_0 (
	.S(\A1[3] ),
	.CO(\CARRYB[5][0] ),
	.CI(\SUMB[4][1] ),
	.B(\CARRYB[4][0] ),
	.A(\ab[5][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_5_1 (
	.S(\SUMB[5][1] ),
	.CO(\CARRYB[5][1] ),
	.CI(\SUMB[4][2] ),
	.B(\CARRYB[4][1] ),
	.A(\ab[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S1_4_0 (
	.S(\A1[2] ),
	.CO(\CARRYB[4][0] ),
	.CI(\SUMB[3][1] ),
	.B(\CARRYB[3][0] ),
	.A(\ab[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_4_1 (
	.S(\SUMB[4][1] ),
	.CO(\CARRYB[4][1] ),
	.CI(\SUMB[3][2] ),
	.B(\CARRYB[3][1] ),
	.A(\ab[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_3_1 (
	.S(\SUMB[3][1] ),
	.CO(\CARRYB[3][1] ),
	.CI(\SUMB[2][2] ),
	.B(\CARRYB[2][1] ),
	.A(\ab[3][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_3_5 (
	.S(\SUMB[3][5] ),
	.CO(\CARRYB[3][5] ),
	.CI(\SUMB[2][6] ),
	.B(\CARRYB[2][5] ),
	.A(\ab[3][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S1_2_0 (
	.S(\A1[0] ),
	.CO(\CARRYB[2][0] ),
	.CI(\SUMB[1][1] ),
	.B(n7),
	.A(\ab[2][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_2_1 (
	.S(\SUMB[2][1] ),
	.CO(\CARRYB[2][1] ),
	.CI(\SUMB[1][2] ),
	.B(n4),
	.A(\ab[2][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_6_5 (
	.S(\SUMB[6][5] ),
	.CO(\CARRYB[6][5] ),
	.CI(\SUMB[5][6] ),
	.B(\CARRYB[5][5] ),
	.A(\ab[6][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S3_5_6 (
	.S(\SUMB[5][6] ),
	.CO(\CARRYB[5][6] ),
	.CI(\ab[4][7] ),
	.B(\CARRYB[4][6] ),
	.A(\ab[5][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_5_5 (
	.S(\SUMB[5][5] ),
	.CO(\CARRYB[5][5] ),
	.CI(\SUMB[4][6] ),
	.B(\CARRYB[4][5] ),
	.A(\ab[5][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S3_4_6 (
	.S(\SUMB[4][6] ),
	.CO(\CARRYB[4][6] ),
	.CI(\ab[3][7] ),
	.B(\CARRYB[3][6] ),
	.A(\ab[4][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_4_5 (
	.S(\SUMB[4][5] ),
	.CO(\CARRYB[4][5] ),
	.CI(\SUMB[3][6] ),
	.B(\CARRYB[3][5] ),
	.A(\ab[4][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S3_3_6 (
	.S(\SUMB[3][6] ),
	.CO(\CARRYB[3][6] ),
	.CI(\ab[2][7] ),
	.B(\CARRYB[2][6] ),
	.A(\ab[3][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S3_2_6 (
	.S(\SUMB[2][6] ),
	.CO(\CARRYB[2][6] ),
	.CI(\ab[1][7] ),
	.B(n9),
	.A(\ab[2][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_2_5 (
	.S(\SUMB[2][5] ),
	.CO(\CARRYB[2][5] ),
	.CI(\SUMB[1][6] ),
	.B(n3),
	.A(\ab[2][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_0 (
	.S(\SUMB[7][0] ),
	.CO(\CARRYB[7][0] ),
	.CI(\SUMB[6][1] ),
	.B(\CARRYB[6][0] ),
	.A(\ab[7][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_1 (
	.S(\SUMB[7][1] ),
	.CO(\CARRYB[7][1] ),
	.CI(\SUMB[6][2] ),
	.B(\CARRYB[6][1] ),
	.A(\ab[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_5 (
	.S(\SUMB[7][5] ),
	.CO(\CARRYB[7][5] ),
	.CI(\SUMB[6][6] ),
	.B(\CARRYB[6][5] ),
	.A(\ab[7][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U2 (
	.Y(n3),
	.B(\ab[1][5] ),
	.A(\ab[0][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U3 (
	.Y(n4),
	.B(\ab[1][1] ),
	.A(\ab[0][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U4 (
	.Y(n5),
	.B(\ab[1][3] ),
	.A(\ab[0][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U5 (
	.Y(n6),
	.B(\ab[1][2] ),
	.A(\ab[0][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U6 (
	.Y(n7),
	.B(\ab[1][0] ),
	.A(\ab[0][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U7 (
	.Y(n8),
	.B(\ab[1][4] ),
	.A(\ab[0][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U8 (
	.Y(n9),
	.B(\ab[1][6] ),
	.A(\ab[0][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U9 (
	.Y(n10),
	.B(\ab[7][7] ),
	.A(\CARRYB[7][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U10 (
	.Y(n23),
	.A(\ab[0][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U11 (
	.Y(n22),
	.A(\ab[0][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U12 (
	.Y(n24),
	.A(\ab[0][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U13 (
	.Y(n11),
	.B(\SUMB[7][1] ),
	.A(\CARRYB[7][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U14 (
	.Y(\A1[11] ),
	.B(\SUMB[7][6] ),
	.A(\CARRYB[7][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U15 (
	.Y(n12),
	.B(\SUMB[7][6] ),
	.A(\CARRYB[7][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U16 (
	.Y(\A1[6] ),
	.B(n17),
	.A(\CARRYB[7][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U17 (
	.Y(n17),
	.A(\SUMB[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U18 (
	.Y(\A1[12] ),
	.B(\ab[7][7] ),
	.A(\CARRYB[7][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U19 (
	.Y(\A1[7] ),
	.B(\SUMB[7][2] ),
	.A(\CARRYB[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U20 (
	.Y(\A1[8] ),
	.B(\SUMB[7][3] ),
	.A(\CARRYB[7][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U21 (
	.Y(\A1[10] ),
	.B(\SUMB[7][5] ),
	.A(\CARRYB[7][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U22 (
	.Y(\A1[9] ),
	.B(\SUMB[7][4] ),
	.A(\CARRYB[7][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U23 (
	.Y(n20),
	.A(\ab[0][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U24 (
	.Y(n21),
	.A(\ab[0][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U25 (
	.Y(n19),
	.A(\ab[0][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U26 (
	.Y(\SUMB[1][6] ),
	.B(n24),
	.A(\ab[1][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U27 (
	.Y(\SUMB[1][2] ),
	.B(n20),
	.A(\ab[1][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U28 (
	.Y(\SUMB[1][1] ),
	.B(n19),
	.A(\ab[1][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U29 (
	.Y(n13),
	.B(\SUMB[7][2] ),
	.A(\CARRYB[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U30 (
	.Y(n14),
	.B(\SUMB[7][3] ),
	.A(\CARRYB[7][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U31 (
	.Y(n15),
	.B(\SUMB[7][4] ),
	.A(\CARRYB[7][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U32 (
	.Y(n16),
	.B(\SUMB[7][5] ),
	.A(\CARRYB[7][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U33 (
	.Y(PRODUCT[1]),
	.B(n18),
	.A(\ab[1][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U34 (
	.Y(n18),
	.A(\ab[0][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U35 (
	.Y(\SUMB[1][5] ),
	.B(n23),
	.A(\ab[1][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U36 (
	.Y(\SUMB[1][4] ),
	.B(n22),
	.A(\ab[1][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U37 (
	.Y(\SUMB[1][3] ),
	.B(n21),
	.A(\ab[1][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U38 (
	.Y(n35),
	.A(B[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U43 (
	.Y(n39),
	.A(B[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U44 (
	.Y(n27),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U47 (
	.Y(n36),
	.A(B[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U48 (
	.Y(n38),
	.A(B[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U49 (
	.Y(n37),
	.A(B[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U50 (
	.Y(n34),
	.A(B[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U51 (
	.Y(n25),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U53 (
	.Y(n40),
	.A(B[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U55 (
	.Y(\ab[7][7] ),
	.B(n177),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U56 (
	.Y(\ab[7][6] ),
	.B(n34),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U57 (
	.Y(\ab[7][5] ),
	.B(n35),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U58 (
	.Y(\ab[7][4] ),
	.B(n36),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U59 (
	.Y(\ab[7][3] ),
	.B(n37),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U60 (
	.Y(\ab[7][2] ),
	.B(n38),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U61 (
	.Y(\ab[7][1] ),
	.B(n39),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U62 (
	.Y(\ab[7][0] ),
	.B(n40),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U63 (
	.Y(\ab[6][7] ),
	.B(n183),
	.A(n177), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U64 (
	.Y(\ab[6][6] ),
	.B(n183),
	.A(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U65 (
	.Y(\ab[6][5] ),
	.B(n183),
	.A(n35), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U66 (
	.Y(\ab[6][4] ),
	.B(n183),
	.A(n36), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U67 (
	.Y(\ab[6][3] ),
	.B(n183),
	.A(n37), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U68 (
	.Y(\ab[6][2] ),
	.B(n183),
	.A(n38), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U69 (
	.Y(\ab[6][1] ),
	.B(n183),
	.A(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U70 (
	.Y(\ab[6][0] ),
	.B(n183),
	.A(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U71 (
	.Y(\ab[5][7] ),
	.B(n27),
	.A(n177), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U72 (
	.Y(\ab[5][6] ),
	.B(n27),
	.A(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U73 (
	.Y(\ab[5][5] ),
	.B(n27),
	.A(n35), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U74 (
	.Y(\ab[5][4] ),
	.B(n27),
	.A(n36), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U75 (
	.Y(\ab[5][3] ),
	.B(n27),
	.A(n37), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U76 (
	.Y(\ab[5][2] ),
	.B(n27),
	.A(n38), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U77 (
	.Y(\ab[5][1] ),
	.B(n27),
	.A(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U78 (
	.Y(\ab[5][0] ),
	.B(n27),
	.A(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U79 (
	.Y(\ab[4][7] ),
	.B(n200),
	.A(n177), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U80 (
	.Y(\ab[4][6] ),
	.B(n200),
	.A(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U81 (
	.Y(\ab[4][5] ),
	.B(n200),
	.A(n35), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U82 (
	.Y(\ab[4][4] ),
	.B(n200),
	.A(n36), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U83 (
	.Y(\ab[4][3] ),
	.B(n200),
	.A(n37), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U84 (
	.Y(\ab[4][2] ),
	.B(n200),
	.A(n38), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U85 (
	.Y(\ab[4][1] ),
	.B(n200),
	.A(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U86 (
	.Y(\ab[4][0] ),
	.B(n200),
	.A(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U87 (
	.Y(\ab[3][7] ),
	.B(n209),
	.A(n177), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U88 (
	.Y(\ab[3][6] ),
	.B(n209),
	.A(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U89 (
	.Y(\ab[3][5] ),
	.B(n209),
	.A(n35), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U90 (
	.Y(\ab[3][4] ),
	.B(n209),
	.A(n36), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U91 (
	.Y(\ab[3][3] ),
	.B(n209),
	.A(n37), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U92 (
	.Y(\ab[3][2] ),
	.B(n209),
	.A(n38), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U93 (
	.Y(\ab[3][1] ),
	.B(n209),
	.A(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U94 (
	.Y(\ab[3][0] ),
	.B(n209),
	.A(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U95 (
	.Y(\ab[2][7] ),
	.B(n229),
	.A(n177), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U96 (
	.Y(\ab[2][6] ),
	.B(n229),
	.A(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U97 (
	.Y(\ab[2][5] ),
	.B(n229),
	.A(n35), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U98 (
	.Y(\ab[2][4] ),
	.B(n229),
	.A(n36), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U99 (
	.Y(\ab[2][3] ),
	.B(n229),
	.A(n37), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U100 (
	.Y(\ab[2][2] ),
	.B(n229),
	.A(n38), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U101 (
	.Y(\ab[2][1] ),
	.B(n229),
	.A(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U102 (
	.Y(\ab[2][0] ),
	.B(n229),
	.A(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U103 (
	.Y(\ab[1][7] ),
	.B(n93),
	.A(n177), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U104 (
	.Y(\ab[1][6] ),
	.B(n93),
	.A(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U105 (
	.Y(\ab[1][5] ),
	.B(n93),
	.A(n35), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U106 (
	.Y(\ab[1][4] ),
	.B(n93),
	.A(n36), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U107 (
	.Y(\ab[1][3] ),
	.B(n93),
	.A(n37), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U108 (
	.Y(\ab[1][2] ),
	.B(n93),
	.A(n38), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U109 (
	.Y(\ab[1][1] ),
	.B(n93),
	.A(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U110 (
	.Y(\ab[1][0] ),
	.B(n93),
	.A(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U111 (
	.Y(\ab[0][7] ),
	.B(n92),
	.A(n177), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U112 (
	.Y(\ab[0][6] ),
	.B(n92),
	.A(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U113 (
	.Y(\ab[0][5] ),
	.B(n92),
	.A(n35), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U114 (
	.Y(\ab[0][4] ),
	.B(n92),
	.A(n36), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U115 (
	.Y(\ab[0][3] ),
	.B(n92),
	.A(n37), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U116 (
	.Y(\ab[0][2] ),
	.B(n92),
	.A(n38), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U117 (
	.Y(\ab[0][1] ),
	.B(n92),
	.A(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U118 (
	.Y(PRODUCT[0]),
	.B(n92),
	.A(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   ALU_DW01_add_1 FS_1 (
	.A({ 1'b0,
		\A1[12] ,
		\A1[11] ,
		\A1[10] ,
		\A1[9] ,
		\A1[8] ,
		\A1[7] ,
		\A1[6] ,
		\SUMB[7][0] ,
		\A1[4] ,
		\A1[3] ,
		\A1[2] ,
		\A1[1] ,
		\A1[0]  }),
	.B({ n10,
		n12,
		n16,
		n15,
		n14,
		n13,
		n11,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0 }),
	.CI(1'b0),
	.SUM({ PRODUCT[15],
		PRODUCT[14],
		PRODUCT[13],
		PRODUCT[12],
		PRODUCT[11],
		PRODUCT[10],
		PRODUCT[9],
		PRODUCT[8],
		PRODUCT[7],
		PRODUCT[6],
		PRODUCT[5],
		PRODUCT[4],
		PRODUCT[3],
		PRODUCT[2] }), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_DW01_add_1 (
	A, 
	B, 
	CI, 
	SUM, 
	CO, 
	VDD, 
	VSS);
   input [13:0] A;
   input [13:0] B;
   input CI;
   output [13:0] SUM;
   output CO;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n1;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;

   // Module instantiations
   AOI21BX2M U2 (
	.Y(n1),
	.B0N(n19),
	.A1(A[12]),
	.A0(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U3 (
	.Y(n15),
	.B(B[7]),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U4 (
	.Y(n9),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U5 (
	.Y(SUM[13]),
	.B(n1),
	.A(B[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U6 (
	.Y(SUM[7]),
	.B(n8),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U7 (
	.Y(n8),
	.A(B[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U8 (
	.Y(SUM[6]),
	.A(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U9 (
	.Y(SUM[0]),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U10 (
	.Y(SUM[1]),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U11 (
	.Y(SUM[2]),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U12 (
	.Y(SUM[3]),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U13 (
	.Y(SUM[4]),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U14 (
	.Y(SUM[5]),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U15 (
	.Y(SUM[9]),
	.B(n11),
	.A(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U16 (
	.Y(n11),
	.B(n13),
	.A(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U17 (
	.Y(SUM[8]),
	.B(n15),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U18 (
	.Y(n14),
	.B(n17),
	.AN(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U19 (
	.Y(n19),
	.B0(B[12]),
	.A1(n18),
	.A0(A[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U20 (
	.Y(SUM[12]),
	.C(n18),
	.B(A[12]),
	.A(B[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21BX1M U21 (
	.Y(n18),
	.B0N(n22),
	.A1(n21),
	.A0(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U22 (
	.Y(SUM[11]),
	.B(n23),
	.A(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U23 (
	.Y(n23),
	.B(n20),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U24 (
	.Y(n20),
	.B(A[11]),
	.A(B[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U25 (
	.Y(n22),
	.B(A[11]),
	.A(B[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OA21X1M U26 (
	.Y(n21),
	.B0(n26),
	.A1(n25),
	.A0(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U27 (
	.Y(SUM[10]),
	.B(n25),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2BB1X1M U28 (
	.Y(n25),
	.B0(n12),
	.A1N(n13),
	.A0N(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U29 (
	.Y(n12),
	.B(A[9]),
	.A(B[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U30 (
	.Y(n13),
	.B(A[9]),
	.A(B[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OA21X1M U31 (
	.Y(n10),
	.B0(n17),
	.A1(n16),
	.A0(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U32 (
	.Y(n17),
	.B(A[8]),
	.A(B[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U33 (
	.Y(n16),
	.B(A[8]),
	.A(B[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U34 (
	.Y(n27),
	.B(n26),
	.AN(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U35 (
	.Y(n26),
	.B(A[10]),
	.A(B[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U36 (
	.Y(n24),
	.B(A[10]),
	.A(B[10]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_DW_div_uns_1 (
	a, 
	b, 
	quotient, 
	remainder, 
	divide_by_0, 
	n200, 
	n209, 
	FE_PT1_n92, 
	FE_PT1_n93, 
	n176, 
	n183, 
	n177, 
	VDD, 
	VSS);
   input [7:0] a;
   input [7:0] b;
   output [7:0] quotient;
   output [7:0] remainder;
   output divide_by_0;
   input n200;
   input n209;
   input FE_PT1_n92;
   input FE_PT1_n93;
   input n176;
   input n183;
   input n177;
   inout VDD;
   inout VSS;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire FE_RN_416_0;
   wire FE_RN_414_0;
   wire FE_RN_413_0;
   wire FE_RN_412_0;
   wire FE_RN_411_0;
   wire FE_RN_410_0;
   wire FE_RN_409_0;
   wire FE_RN_408_0;
   wire FE_RN_407_0;
   wire FE_RN_406_0;
   wire FE_RN_403_0;
   wire FE_RN_402_0;
   wire FE_RN_338_0;
   wire FE_RN_337_0;
   wire FE_RN_336_0;
   wire FE_RN_335_0;
   wire FE_RN_334_0;
   wire FE_RN_333_0;
   wire FE_RN_332_0;
   wire FE_RN_331_0;
   wire FE_RN_330_0;
   wire FE_RN_329_0;
   wire FE_RN_328_0;
   wire FE_RN_327_0;
   wire FE_RN_326_0;
   wire FE_RN_325_0;
   wire FE_RN_324_0;
   wire FE_RN_323_0;
   wire FE_RN_322_0;
   wire FE_RN_321_0;
   wire FE_RN_320_0;
   wire FE_RN_316_0;
   wire FE_RN_315_0;
   wire FE_RN_314_0;
   wire FE_RN_313_0;
   wire FE_RN_312_0;
   wire FE_RN_311_0;
   wire FE_RN_310_0;
   wire FE_RN_309_0;
   wire FE_RN_308_0;
   wire FE_RN_307_0;
   wire FE_RN_306_0;
   wire FE_RN_304_0;
   wire FE_RN_303_0;
   wire FE_RN_302_0;
   wire FE_RN_299_0;
   wire FE_RN_298_0;
   wire FE_RN_297_0;
   wire FE_RN_295_0;
   wire FE_RN_294_0;
   wire FE_RN_293_0;
   wire FE_RN_292_0;
   wire FE_RN_291_0;
   wire FE_RN_290_0;
   wire FE_RN_289_0;
   wire FE_RN_288_0;
   wire FE_RN_287_0;
   wire FE_RN_207_0;
   wire FE_RN_206_0;
   wire FE_RN_205_0;
   wire FE_RN_204_0;
   wire FE_RN_203_0;
   wire FE_RN_202_0;
   wire FE_RN_201_0;
   wire FE_RN_200_0;
   wire FE_RN_199_0;
   wire FE_RN_198_0;
   wire FE_RN_197_0;
   wire FE_RN_196_0;
   wire FE_RN_195_0;
   wire FE_RN_194_0;
   wire FE_RN_193_0;
   wire FE_RN_192_0;
   wire FE_RN_191_0;
   wire FE_RN_190_0;
   wire FE_RN_189_0;
   wire FE_RN_188_0;
   wire FE_RN_187_0;
   wire FE_RN_109_0;
   wire FE_RN_108_0;
   wire FE_RN_106_0;
   wire FE_RN_105_0;
   wire FE_RN_104_0;
   wire FE_RN_103_0;
   wire FE_RN_71_0;
   wire FE_RN_70_0;
   wire FE_RN_69_0;
   wire FE_RN_68_0;
   wire FE_RN_67_0;
   wire FE_RN_66_0;
   wire FE_RN_65_0;
   wire FE_RN_64_0;
   wire FE_RN_63_0;
   wire FE_RN_62_0;
   wire FE_RN_61_0;
   wire FE_RN_60_0;
   wire FE_RN_59_0;
   wire FE_RN_58_0;
   wire FE_RN_57_0;
   wire FE_RN_56_0;
   wire FE_RN_55_0;
   wire FE_RN_54_0;
   wire FE_RN_53_0;
   wire FE_RN_52_0;
   wire FE_RN_51_0;
   wire FE_RN_50_0;
   wire FE_RN_49_0;
   wire FE_RN_47_0;
   wire FE_RN_46_0;
   wire FE_RN_45_0;
   wire FE_OFN13_N127;
   wire \u_div/SumTmp[1][1] ;
   wire \u_div/SumTmp[1][2] ;
   wire \u_div/SumTmp[1][3] ;
   wire \u_div/SumTmp[1][4] ;
   wire \u_div/SumTmp[1][5] ;
   wire \u_div/SumTmp[1][6] ;
   wire \u_div/SumTmp[2][0] ;
   wire \u_div/SumTmp[2][1] ;
   wire \u_div/SumTmp[2][2] ;
   wire \u_div/SumTmp[2][3] ;
   wire \u_div/SumTmp[2][4] ;
   wire \u_div/SumTmp[2][5] ;
   wire \u_div/SumTmp[3][0] ;
   wire \u_div/SumTmp[3][1] ;
   wire \u_div/SumTmp[3][2] ;
   wire \u_div/SumTmp[3][3] ;
   wire \u_div/SumTmp[3][4] ;
   wire \u_div/SumTmp[4][0] ;
   wire \u_div/SumTmp[4][1] ;
   wire \u_div/SumTmp[4][2] ;
   wire \u_div/SumTmp[4][3] ;
   wire \u_div/SumTmp[5][0] ;
   wire \u_div/SumTmp[5][1] ;
   wire \u_div/SumTmp[5][2] ;
   wire \u_div/SumTmp[6][0] ;
   wire \u_div/SumTmp[6][1] ;
   wire \u_div/CryTmp[0][1] ;
   wire \u_div/CryTmp[0][2] ;
   wire \u_div/CryTmp[0][3] ;
   wire \u_div/CryTmp[0][4] ;
   wire \u_div/CryTmp[0][5] ;
   wire \u_div/CryTmp[0][6] ;
   wire \u_div/CryTmp[0][7] ;
   wire \u_div/CryTmp[1][1] ;
   wire \u_div/CryTmp[1][2] ;
   wire \u_div/CryTmp[1][3] ;
   wire \u_div/CryTmp[1][4] ;
   wire \u_div/CryTmp[1][5] ;
   wire \u_div/CryTmp[1][6] ;
   wire \u_div/CryTmp[1][7] ;
   wire \u_div/CryTmp[2][1] ;
   wire \u_div/CryTmp[2][3] ;
   wire \u_div/CryTmp[2][4] ;
   wire \u_div/CryTmp[2][5] ;
   wire \u_div/CryTmp[3][1] ;
   wire \u_div/CryTmp[3][2] ;
   wire \u_div/CryTmp[3][3] ;
   wire \u_div/CryTmp[4][1] ;
   wire \u_div/CryTmp[4][2] ;
   wire \u_div/CryTmp[4][3] ;
   wire \u_div/CryTmp[5][1] ;
   wire \u_div/CryTmp[5][2] ;
   wire \u_div/CryTmp[6][1] ;
   wire \u_div/CryTmp[6][2] ;
   wire \u_div/CryTmp[7][1] ;
   wire \u_div/PartRem[1][1] ;
   wire \u_div/PartRem[1][2] ;
   wire \u_div/PartRem[1][3] ;
   wire \u_div/PartRem[1][4] ;
   wire \u_div/PartRem[1][5] ;
   wire \u_div/PartRem[1][6] ;
   wire \u_div/PartRem[1][7] ;
   wire \u_div/PartRem[2][1] ;
   wire \u_div/PartRem[2][2] ;
   wire \u_div/PartRem[2][3] ;
   wire \u_div/PartRem[2][4] ;
   wire \u_div/PartRem[2][5] ;
   wire \u_div/PartRem[2][6] ;
   wire \u_div/PartRem[4][1] ;
   wire \u_div/PartRem[5][1] ;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n21;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n33;
   wire n34;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n71;
   wire n73;
   wire n74;
   wire n75;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire [7:0] \u_div/BInv ;

   // Module instantiations
   CLKAND2X6M FE_RC_543_0 (
	.Y(n68),
	.B(FE_RN_62_0),
	.A(FE_RN_56_0), 
	.VDD(VDD), 
	.VSS(VSS));
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_542_0 (
	.Y(FE_RN_416_0),
	.A(FE_RN_402_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21BX4M FE_RC_540_0 (
	.Y(n82),
	.B0N(FE_RN_410_0),
	.A1(FE_RN_416_0),
	.A0(\u_div/CryTmp[2][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_539_0 (
	.Y(FE_RN_414_0),
	.A(n81), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX2M FE_RC_538_0 (
	.Y(FE_RN_413_0),
	.C(FE_RN_411_0),
	.B(FE_RN_414_0),
	.AN(FE_RN_402_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_537_0 (
	.Y(FE_RN_412_0),
	.A(\u_div/BInv [5]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M FE_RC_536_0 (
	.Y(FE_RN_411_0),
	.B(FE_RN_412_0),
	.AN(n45), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_535_0 (
	.Y(FE_RN_410_0),
	.A(FE_RN_411_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M FE_RC_534_0 (
	.Y(FE_RN_409_0),
	.B(n81),
	.A(FE_RN_410_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X4M FE_RC_533_0 (
	.Y(FE_RN_408_0),
	.B(\u_div/CryTmp[2][5] ),
	.A(FE_RN_409_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_532_0 (
	.Y(n80),
	.B(FE_RN_413_0),
	.A(FE_RN_408_0), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M FE_RC_531_0 (
	.Y(FE_RN_407_0),
	.B(\u_div/BInv [5]),
	.A(n45), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_530_0 (
	.Y(FE_RN_406_0),
	.A(n45), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M FE_RC_527_0 (
	.Y(FE_RN_403_0),
	.B0(FE_RN_416_0),
	.A1(FE_RN_412_0),
	.A0(FE_RN_406_0), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M FE_RC_526_0 (
	.Y(\u_div/SumTmp[2][5] ),
	.S0(\u_div/CryTmp[2][5] ),
	.B(FE_RN_403_0),
	.A(FE_RN_407_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_525_0 (
	.Y(FE_RN_402_0),
	.B(\u_div/BInv [5]),
	.A(n45), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_447_0 (
	.Y(FE_RN_338_0),
	.A(FE_RN_291_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX2M FE_RC_446_0 (
	.Y(n78),
	.C(FE_RN_201_0),
	.B(FE_RN_187_0),
	.AN(FE_RN_338_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_445_0 (
	.Y(FE_RN_337_0),
	.A(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M FE_RC_444_0 (
	.Y(FE_RN_336_0),
	.B(FE_RN_337_0),
	.AN(FE_RN_289_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M FE_RC_443_0 (
	.Y(n21),
	.B(FE_RN_336_0),
	.AN(FE_RN_299_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_442_0 (
	.Y(FE_RN_335_0),
	.A(\u_div/CryTmp[2][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M FE_RC_441_0 (
	.Y(FE_RN_334_0),
	.C(FE_RN_335_0),
	.B(n209),
	.A(FE_RN_323_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_440_0 (
	.Y(FE_RN_333_0),
	.A(n209), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX2M FE_RC_439_0 (
	.Y(FE_RN_332_0),
	.C(FE_RN_295_0),
	.B(FE_RN_333_0),
	.AN(FE_RN_323_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_438_0 (
	.Y(FE_RN_331_0),
	.B(FE_RN_334_0),
	.A(FE_RN_332_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_437_0 (
	.Y(FE_RN_330_0),
	.A(FE_RN_316_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M FE_RC_436_0 (
	.Y(FE_RN_329_0),
	.B(FE_RN_289_0),
	.A(FE_RN_330_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_435_0 (
	.Y(FE_RN_328_0),
	.A(\u_div/BInv [1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X1M FE_RC_434_0 (
	.Y(FE_RN_327_0),
	.C(FE_RN_328_0),
	.B(n209),
	.A(FE_RN_289_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_433_0 (
	.Y(FE_RN_326_0),
	.B(FE_RN_295_0),
	.A(FE_RN_327_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M FE_RC_432_0 (
	.Y(FE_RN_325_0),
	.B0(FE_RN_326_0),
	.A1(n23),
	.A0(FE_RN_329_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_431_0 (
	.Y(FE_RN_324_0),
	.A(FE_RN_288_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M FE_RC_430_0 (
	.Y(FE_RN_323_0),
	.B(\u_div/BInv [2]),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M FE_RC_429_0 (
	.Y(FE_RN_322_0),
	.B0(FE_RN_323_0),
	.A1(FE_RN_316_0),
	.A0(FE_RN_324_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2B1X1M FE_RC_428_0 (
	.Y(FE_RN_321_0),
	.B0(FE_RN_322_0),
	.A1N(FE_RN_325_0),
	.A0(FE_RN_323_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M FE_RC_427_0 (
	.Y(\u_div/SumTmp[2][2] ),
	.B0(FE_RN_321_0),
	.A1N(FE_RN_331_0),
	.A0N(FE_RN_289_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_426_0 (
	.Y(FE_RN_320_0),
	.B(FE_RN_295_0),
	.A(FE_RN_316_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_422_0 (
	.Y(FE_RN_316_0),
	.B(\u_div/CryTmp[2][1] ),
	.A(\u_div/BInv [1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B1X2M FE_RC_421_0 (
	.Y(FE_RN_315_0),
	.B0(FE_RN_316_0),
	.A1N(FE_RN_328_0),
	.A0(\u_div/CryTmp[2][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M FE_RC_420_0 (
	.Y(FE_RN_314_0),
	.B(FE_RN_337_0),
	.A(FE_RN_315_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M FE_RC_419_0 (
	.Y(FE_RN_313_0),
	.B0(FE_RN_314_0),
	.A1(FE_RN_337_0),
	.A0(FE_RN_320_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_418_0 (
	.Y(FE_RN_312_0),
	.B(\u_div/BInv [1]),
	.A(n209), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M FE_RC_417_0 (
	.Y(FE_RN_311_0),
	.B0(FE_RN_312_0),
	.A1(\u_div/BInv [1]),
	.A0(n209), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_416_0 (
	.Y(FE_RN_310_0),
	.A(FE_RN_311_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_415_0 (
	.Y(FE_RN_309_0),
	.A(\u_div/CryTmp[2][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M FE_RC_414_0 (
	.Y(FE_RN_308_0),
	.B(\u_div/BInv [1]),
	.A(n209), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M FE_RC_413_0 (
	.Y(FE_RN_307_0),
	.B(n209),
	.A(FE_RN_295_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM FE_RC_412_0 (
	.Y(FE_RN_306_0),
	.C0(FE_RN_307_0),
	.B1(FE_RN_308_0),
	.B0(FE_RN_309_0),
	.A1(\u_div/CryTmp[2][1] ),
	.A0(FE_RN_310_0), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M FE_RC_411_0 (
	.Y(\u_div/SumTmp[2][1] ),
	.S0(FE_RN_289_0),
	.B(FE_RN_306_0),
	.A(FE_RN_313_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX2M FE_RC_409_0 (
	.Y(FE_RN_304_0),
	.C(FE_RN_316_0),
	.B(FE_RN_298_0),
	.AN(FE_RN_288_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_408_0 (
	.Y(FE_RN_303_0),
	.B(\u_div/BInv [2]),
	.A(FE_RN_304_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_407_0 (
	.Y(FE_RN_302_0),
	.A(\u_div/BInv [2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M FE_RC_404_0 (
	.Y(FE_RN_299_0),
	.B(FE_RN_333_0),
	.A(FE_RN_289_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_403_0 (
	.Y(FE_RN_298_0),
	.B(FE_RN_295_0),
	.A(FE_RN_299_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X4M FE_RC_402_0 (
	.Y(FE_RN_297_0),
	.C(FE_RN_302_0),
	.B(FE_RN_316_0),
	.A(FE_RN_298_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M FE_RC_400_0 (
	.Y(FE_RN_295_0),
	.B(FE_RN_328_0),
	.AN(\u_div/CryTmp[2][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_399_0 (
	.Y(FE_RN_294_0),
	.A(FE_RN_295_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_398_0 (
	.Y(FE_RN_293_0),
	.A(n77), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_397_0 (
	.Y(FE_RN_292_0),
	.A(FE_RN_190_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_396_0 (
	.Y(FE_RN_291_0),
	.B(FE_RN_188_0),
	.A(FE_RN_292_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M FE_RC_395_0 (
	.Y(FE_RN_290_0),
	.B(FE_RN_201_0),
	.A(FE_RN_291_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X4M FE_RC_394_0 (
	.Y(FE_RN_289_0),
	.C(FE_RN_293_0),
	.B(FE_RN_187_0),
	.A(FE_RN_290_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X4M FE_RC_393_0 (
	.Y(FE_RN_288_0),
	.C(n23),
	.B(FE_RN_294_0),
	.A(FE_RN_289_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X4M FE_RC_392_0 (
	.Y(FE_RN_287_0),
	.B0(n1),
	.A1(FE_RN_288_0),
	.A0(FE_RN_297_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_391_0 (
	.Y(\u_div/CryTmp[2][3] ),
	.B(FE_RN_303_0),
	.A(FE_RN_287_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX2M FE_RC_300_0 (
	.Y(FE_RN_207_0),
	.C(FE_RN_189_0),
	.B(FE_RN_205_0),
	.AN(\u_div/CryTmp[3][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_299_0 (
	.Y(FE_RN_206_0),
	.A(FE_RN_190_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M FE_RC_298_0 (
	.Y(FE_RN_205_0),
	.B(\u_div/BInv [4]),
	.A(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_297_0 (
	.Y(FE_RN_204_0),
	.B(FE_RN_206_0),
	.A(FE_RN_205_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_296_0 (
	.Y(FE_RN_203_0),
	.A(\u_div/BInv [4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_295_0 (
	.Y(FE_RN_202_0),
	.A(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_294_0 (
	.Y(FE_RN_201_0),
	.B(FE_RN_203_0),
	.A(FE_RN_202_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_293_0 (
	.Y(FE_RN_200_0),
	.B(FE_RN_188_0),
	.A(FE_RN_201_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_292_0 (
	.Y(FE_RN_199_0),
	.B(\u_div/CryTmp[3][3] ),
	.A(FE_RN_190_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_291_0 (
	.Y(FE_RN_198_0),
	.B(FE_RN_189_0),
	.A(FE_RN_199_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_290_0 (
	.Y(FE_RN_197_0),
	.B(FE_RN_200_0),
	.A(FE_RN_198_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M FE_RC_289_0 (
	.Y(\u_div/SumTmp[3][4] ),
	.C(FE_RN_207_0),
	.B(FE_RN_204_0),
	.A(FE_RN_197_0), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR2X2M FE_RC_288_0 (
	.Y(FE_RN_196_0),
	.B(\u_div/BInv [3]),
	.A(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M FE_RC_287_0 (
	.Y(FE_RN_195_0),
	.B(FE_RN_196_0),
	.AN(\u_div/CryTmp[3][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_286_0 (
	.Y(FE_RN_194_0),
	.B(FE_RN_189_0),
	.A(FE_RN_190_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_285_0 (
	.Y(FE_RN_193_0),
	.B(\u_div/CryTmp[3][3] ),
	.A(FE_RN_194_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_284_0 (
	.Y(\u_div/SumTmp[3][3] ),
	.B(FE_RN_195_0),
	.A(FE_RN_193_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_283_0 (
	.Y(FE_RN_192_0),
	.A(\u_div/BInv [3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_282_0 (
	.Y(FE_RN_191_0),
	.A(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_281_0 (
	.Y(FE_RN_190_0),
	.B(FE_RN_192_0),
	.A(FE_RN_191_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_280_0 (
	.Y(FE_RN_189_0),
	.B(\u_div/BInv [3]),
	.A(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_279_0 (
	.Y(FE_RN_188_0),
	.B(\u_div/BInv [4]),
	.A(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX4M FE_RC_278_0 (
	.Y(FE_RN_187_0),
	.C(FE_RN_188_0),
	.B(FE_RN_189_0),
	.AN(\u_div/CryTmp[3][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_183_0 (
	.Y(n74),
	.A(FE_RN_104_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_182_0 (
	.Y(FE_RN_109_0),
	.A(n73), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_181_0 (
	.Y(FE_RN_108_0),
	.A(n43), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_179_0 (
	.Y(FE_RN_106_0),
	.B(FE_RN_108_0),
	.A(FE_RN_192_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_178_0 (
	.Y(FE_RN_105_0),
	.B(\u_div/CryTmp[4][3] ),
	.A(FE_RN_106_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_177_0 (
	.Y(FE_RN_104_0),
	.B(n12),
	.A(FE_RN_105_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_176_0 (
	.Y(FE_RN_103_0),
	.B(FE_RN_109_0),
	.A(FE_RN_104_0), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X3M FE_RC_175_0 (
	.Y(\u_div/PartRem[4][1] ),
	.S0(FE_RN_103_0),
	.B(n200),
	.A(n71), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_121_0 (
	.Y(FE_RN_71_0),
	.A(FE_RN_57_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_120_0 (
	.Y(n36),
	.B(FE_RN_59_0),
	.A(FE_RN_71_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_119_0 (
	.Y(FE_RN_70_0),
	.A(\u_div/BInv [2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_118_0 (
	.Y(FE_RN_69_0),
	.A(\u_div/BInv [2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M FE_RC_117_0 (
	.Y(FE_RN_68_0),
	.B1(FE_RN_69_0),
	.B0(\u_div/SumTmp[6][1] ),
	.A1N(\u_div/SumTmp[6][1] ),
	.A0N(FE_RN_70_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_116_0 (
	.Y(FE_RN_67_0),
	.A(\u_div/BInv [2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_115_0 (
	.Y(FE_RN_66_0),
	.A(\u_div/BInv [2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M FE_RC_114_0 (
	.Y(FE_RN_65_0),
	.B1(FE_RN_66_0),
	.B0(n47),
	.A1N(n47),
	.A0N(FE_RN_67_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_113_0 (
	.Y(FE_RN_64_0),
	.A(quotient[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M FE_RC_112_0 (
	.Y(FE_RN_63_0),
	.S0(FE_RN_64_0),
	.B(FE_RN_65_0),
	.A(FE_RN_68_0), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M FE_RC_111_0 (
	.Y(\u_div/SumTmp[5][2] ),
	.B(\u_div/CryTmp[5][2] ),
	.A(FE_RN_63_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M FE_RC_110_0 (
	.Y(FE_RN_62_0),
	.B0(\u_div/BInv [2]),
	.A1(FE_RN_57_0),
	.A0(FE_RN_60_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_109_0 (
	.Y(FE_RN_61_0),
	.A(\u_div/BInv [2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M FE_RC_108_0 (
	.Y(FE_RN_60_0),
	.B(quotient[6]),
	.AN(n47), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_107_0 (
	.Y(FE_RN_59_0),
	.A(FE_RN_60_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_106_0 (
	.Y(FE_RN_58_0),
	.B(FE_RN_61_0),
	.A(FE_RN_59_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M FE_RC_105_0 (
	.Y(FE_RN_57_0),
	.B(quotient[6]),
	.A(\u_div/SumTmp[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M FE_RC_104_0 (
	.Y(FE_RN_56_0),
	.B0(\u_div/CryTmp[5][2] ),
	.A1(FE_RN_57_0),
	.A0(FE_RN_58_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_102_0 (
	.Y(quotient[6]),
	.A(n87), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_101_0 (
	.Y(n34),
	.B(FE_RN_50_0),
	.A(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M FE_RC_100_0 (
	.Y(FE_RN_55_0),
	.B(FE_RN_45_0),
	.AN(FE_RN_47_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_99_0 (
	.Y(FE_RN_54_0),
	.A(FE_RN_45_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M FE_RC_98_0 (
	.Y(FE_RN_53_0),
	.B0(FE_RN_54_0),
	.A1(\u_div/CryTmp[5][1] ),
	.A0(\u_div/BInv [1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_97_0 (
	.Y(FE_RN_52_0),
	.A(FE_RN_53_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_96_0 (
	.Y(FE_RN_51_0),
	.B(FE_RN_52_0),
	.A(FE_RN_49_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M FE_RC_95_0 (
	.Y(\u_div/SumTmp[5][1] ),
	.B0(FE_RN_51_0),
	.A1(FE_RN_49_0),
	.A0(FE_RN_55_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M FE_RC_94_0 (
	.Y(FE_RN_50_0),
	.B(n62),
	.AN(n87), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_93_0 (
	.Y(FE_RN_49_0),
	.B(n33),
	.A(FE_RN_50_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M FE_RC_91_0 (
	.Y(FE_RN_47_0),
	.B(FE_RN_328_0),
	.AN(\u_div/CryTmp[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_90_0 (
	.Y(FE_RN_46_0),
	.A(FE_RN_47_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M FE_RC_89_0 (
	.Y(FE_RN_45_0),
	.B(\u_div/CryTmp[5][1] ),
	.A(\u_div/BInv [1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21BX4M FE_RC_88_0 (
	.Y(\u_div/CryTmp[5][2] ),
	.B0N(FE_RN_45_0),
	.A1(FE_RN_46_0),
	.A0(FE_RN_49_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M FE_RC_8_0 (
	.Y(\u_div/BInv [7]),
	.A(b[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_5_0 (
	.Y(n81),
	.B(\u_div/BInv [6]),
	.A(n177), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X6M FE_RC_4_0 (
	.Y(n91),
	.B(b[7]),
	.A(b[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX8M FE_OFC13_N127 (
	.Y(quotient[3]),
	.A(FE_OFN13_N127), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX4M \u_div/u_fa_PartRem_0_2_4  (
	.S(\u_div/SumTmp[2][4] ),
	.CO(\u_div/CryTmp[2][5] ),
	.CI(\u_div/CryTmp[2][4] ),
	.B(\u_div/BInv [4]),
	.A(n44), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX4M \u_div/u_fa_PartRem_0_2_3  (
	.S(\u_div/SumTmp[2][3] ),
	.CO(\u_div/CryTmp[2][4] ),
	.CI(\u_div/CryTmp[2][3] ),
	.B(\u_div/BInv [3]),
	.A(n42), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX4M \u_div/u_fa_PartRem_0_0_2  (
	.CO(\u_div/CryTmp[0][3] ),
	.CI(\u_div/CryTmp[0][2] ),
	.B(\u_div/BInv [2]),
	.A(\u_div/PartRem[1][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX4M \u_div/u_fa_PartRem_0_0_3  (
	.CO(\u_div/CryTmp[0][4] ),
	.CI(\u_div/CryTmp[0][3] ),
	.B(\u_div/BInv [3]),
	.A(\u_div/PartRem[1][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX4M \u_div/u_fa_PartRem_0_0_1  (
	.CO(\u_div/CryTmp[0][2] ),
	.CI(\u_div/PartRem[1][1] ),
	.B(\u_div/BInv [1]),
	.A(\u_div/CryTmp[0][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX2M \u_div/u_fa_PartRem_0_3_1  (
	.S(\u_div/SumTmp[3][1] ),
	.CO(\u_div/CryTmp[3][2] ),
	.CI(\u_div/CryTmp[3][1] ),
	.B(\u_div/BInv [1]),
	.A(\u_div/PartRem[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX4M \u_div/u_fa_PartRem_0_0_5  (
	.CO(\u_div/CryTmp[0][6] ),
	.CI(\u_div/CryTmp[0][5] ),
	.B(\u_div/BInv [5]),
	.A(\u_div/PartRem[1][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX4M \u_div/u_fa_PartRem_0_0_6  (
	.CO(\u_div/CryTmp[0][7] ),
	.CI(\u_div/CryTmp[0][6] ),
	.B(\u_div/BInv [6]),
	.A(\u_div/PartRem[1][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX4M \u_div/u_fa_PartRem_0_0_4  (
	.CO(\u_div/CryTmp[0][5] ),
	.CI(\u_div/CryTmp[0][4] ),
	.B(\u_div/BInv [4]),
	.A(\u_div/PartRem[1][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX4M \u_div/u_fa_PartRem_0_3_2  (
	.S(\u_div/SumTmp[3][2] ),
	.CO(\u_div/CryTmp[3][3] ),
	.CI(\u_div/CryTmp[3][2] ),
	.B(\u_div/BInv [2]),
	.A(n41), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX4M \u_div/u_fa_PartRem_0_1_1  (
	.S(\u_div/SumTmp[1][1] ),
	.CO(\u_div/CryTmp[1][2] ),
	.CI(\u_div/CryTmp[1][1] ),
	.B(\u_div/BInv [1]),
	.A(\u_div/PartRem[2][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX4M \u_div/u_fa_PartRem_0_1_2  (
	.S(\u_div/SumTmp[1][2] ),
	.CO(\u_div/CryTmp[1][3] ),
	.CI(\u_div/CryTmp[1][2] ),
	.B(\u_div/BInv [2]),
	.A(\u_div/PartRem[2][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX4M \u_div/u_fa_PartRem_0_1_5  (
	.S(\u_div/SumTmp[1][5] ),
	.CO(\u_div/CryTmp[1][6] ),
	.CI(\u_div/CryTmp[1][5] ),
	.B(\u_div/BInv [5]),
	.A(\u_div/PartRem[2][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX4M \u_div/u_fa_PartRem_0_1_3  (
	.S(\u_div/SumTmp[1][3] ),
	.CO(\u_div/CryTmp[1][4] ),
	.CI(\u_div/CryTmp[1][3] ),
	.B(\u_div/BInv [3]),
	.A(\u_div/PartRem[2][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX4M \u_div/u_fa_PartRem_0_1_4  (
	.S(\u_div/SumTmp[1][4] ),
	.CO(\u_div/CryTmp[1][5] ),
	.CI(\u_div/CryTmp[1][4] ),
	.B(\u_div/BInv [4]),
	.A(\u_div/PartRem[2][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX4M \u_div/u_fa_PartRem_0_1_6  (
	.S(\u_div/SumTmp[1][6] ),
	.CO(\u_div/CryTmp[1][7] ),
	.CI(\u_div/CryTmp[1][6] ),
	.B(\u_div/BInv [6]),
	.A(\u_div/PartRem[2][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR2XLM U2 (
	.Y(n5),
	.B(\u_div/BInv [2]),
	.A(n37), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2XLM U3 (
	.Y(n40),
	.S0(n27),
	.B(\u_div/SumTmp[4][2] ),
	.A(n37), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X2M U4 (
	.Y(n37),
	.S0(quotient[5]),
	.B(n38),
	.A(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U7 (
	.Y(n2),
	.B(\u_div/BInv [1]),
	.A(\u_div/PartRem[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U11 (
	.Y(\u_div/CryTmp[7][1] ),
	.B(a[7]),
	.A(\u_div/BInv [0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U12 (
	.Y(n84),
	.B(n86),
	.A(n85), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M U13 (
	.Y(n73),
	.B(n91),
	.A(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U15 (
	.Y(n24),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M U16 (
	.Y(n67),
	.B(\u_div/BInv [3]),
	.A(n89), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX4M U17 (
	.Y(n89),
	.A(n73), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U20 (
	.Y(n8),
	.B(\u_div/CryTmp[4][2] ),
	.A(\u_div/BInv [2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U21 (
	.Y(\u_div/CryTmp[4][2] ),
	.C(n4),
	.B(n3),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X4M U22 (
	.Y(n1),
	.S0(quotient[3]),
	.B(\u_div/SumTmp[3][1] ),
	.A(\u_div/PartRem[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX4M U23 (
	.Y(quotient[2]),
	.A(n92), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX4M U24 (
	.Y(quotient[1]),
	.A(n93), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X6M U25 (
	.Y(\u_div/PartRem[1][1] ),
	.S0(n83),
	.B(n50),
	.A(FE_PT1_n93), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX8M U26 (
	.Y(n83),
	.B(b[7]),
	.AN(\u_div/CryTmp[1][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X1M U27 (
	.Y(n43),
	.S0(quotient[5]),
	.B(\u_div/SumTmp[5][2] ),
	.A(n36), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X3M U28 (
	.Y(n57),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][1] ),
	.A(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U31 (
	.Y(\u_div/PartRem[1][3] ),
	.S0(quotient[1]),
	.B(n75),
	.A(n57), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX4M U32 (
	.Y(n86),
	.A(n67), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U33 (
	.Y(n90),
	.B(b[4]),
	.A(b[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX6M U34 (
	.Y(\u_div/BInv [3]),
	.A(b[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX4M U35 (
	.Y(\u_div/BInv [1]),
	.A(b[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U36 (
	.Y(quotient[5]),
	.A(n88), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U37 (
	.Y(quotient[7]),
	.A(n84), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U39 (
	.Y(n3),
	.B(\u_div/CryTmp[4][1] ),
	.A(\u_div/PartRem[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X3M U42 (
	.Y(\u_div/PartRem[5][1] ),
	.S0(n66),
	.B(n65),
	.A(n64), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3BX4M U43 (
	.Y(n85),
	.C(b[1]),
	.B(b[2]),
	.AN(\u_div/CryTmp[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX8M U45 (
	.Y(\u_div/BInv [0]),
	.A(b[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U46 (
	.Y(\u_div/SumTmp[4][1] ),
	.C(\u_div/CryTmp[4][1] ),
	.B(\u_div/BInv [1]),
	.A(\u_div/PartRem[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U47 (
	.Y(n4),
	.B(\u_div/CryTmp[4][1] ),
	.A(\u_div/BInv [1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U48 (
	.Y(\u_div/SumTmp[4][2] ),
	.B(\u_div/CryTmp[4][2] ),
	.A(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U49 (
	.Y(n6),
	.B(\u_div/BInv [2]),
	.A(n37), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U50 (
	.Y(n7),
	.B(\u_div/CryTmp[4][2] ),
	.A(n37), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U51 (
	.Y(\u_div/CryTmp[4][3] ),
	.C(n8),
	.B(n7),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR2XLM U52 (
	.Y(n9),
	.B(n43),
	.A(\u_div/BInv [3]), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR2XLM U53 (
	.Y(\u_div/SumTmp[4][3] ),
	.B(\u_div/CryTmp[4][3] ),
	.A(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U54 (
	.Y(n12),
	.B(\u_div/BInv [3]),
	.A(n43), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR2XLM U56 (
	.Y(n13),
	.B(\u_div/BInv [1]),
	.A(\u_div/CryTmp[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR2X1M U57 (
	.Y(\u_div/SumTmp[6][1] ),
	.B(n47),
	.A(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U58 (
	.Y(n14),
	.B(\u_div/BInv [1]),
	.A(n47), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U59 (
	.Y(n15),
	.B(\u_div/CryTmp[6][1] ),
	.A(n47), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U60 (
	.Y(n16),
	.B(\u_div/CryTmp[6][1] ),
	.A(\u_div/BInv [1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U61 (
	.Y(\u_div/CryTmp[6][2] ),
	.C(n14),
	.B(n15),
	.A(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX4M U62 (
	.Y(n47),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U63 (
	.Y(n87),
	.B(n46),
	.A(\u_div/CryTmp[6][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U64 (
	.Y(n17),
	.B(\u_div/PartRem[1][7] ),
	.A(\u_div/CryTmp[0][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U65 (
	.Y(n18),
	.B(\u_div/BInv [7]),
	.A(\u_div/CryTmp[0][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2XLM U66 (
	.Y(n19),
	.B(\u_div/BInv [7]),
	.A(\u_div/PartRem[1][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U67 (
	.Y(quotient[0]),
	.C(n17),
	.B(n18),
	.A(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2XLM U68 (
	.Y(n28),
	.B(n84),
	.A(n48), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X4M U72 (
	.Y(n27),
	.B(n73),
	.A(n74), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U73 (
	.Y(FE_OFN13_N127),
	.B(n77),
	.A(n78), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X4M U74 (
	.Y(n66),
	.B(n67),
	.A(n68), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX4M U75 (
	.Y(\u_div/PartRem[2][1] ),
	.A(n58), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX4M U76 (
	.Y(\u_div/PartRem[2][2] ),
	.A(n57), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X1M U77 (
	.Y(n33),
	.B(n87),
	.A(n61), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U78 (
	.Y(n93),
	.B(\u_div/CryTmp[1][7] ),
	.AN(b[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U79 (
	.Y(n41),
	.B(n26),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U80 (
	.Y(n23),
	.A(\u_div/SumTmp[3][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U82 (
	.Y(quotient[4]),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U83 (
	.Y(n65),
	.A(\u_div/SumTmp[5][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U84 (
	.Y(\u_div/BInv [2]),
	.A(b[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U85 (
	.Y(n42),
	.S0(quotient[3]),
	.B(\u_div/SumTmp[3][2] ),
	.A(n41), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U87 (
	.Y(n62),
	.A(\u_div/SumTmp[6][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U88 (
	.Y(n92),
	.B(n91),
	.AN(n82), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U89 (
	.Y(\u_div/CryTmp[1][1] ),
	.B(FE_PT1_n93),
	.AN(\u_div/BInv [0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U90 (
	.Y(n61),
	.A(a[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2XLM U91 (
	.Y(n25),
	.B(n24),
	.A(\u_div/PartRem[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2XLM U92 (
	.Y(n26),
	.B(n27),
	.A(\u_div/SumTmp[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U93 (
	.Y(n88),
	.B(n86),
	.AN(n68), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U94 (
	.Y(n79),
	.A(\u_div/SumTmp[1][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U95 (
	.Y(n38),
	.A(\u_div/SumTmp[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X4M U96 (
	.Y(n58),
	.S0(n80),
	.B(\u_div/SumTmp[2][0] ),
	.A(a[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U97 (
	.Y(\u_div/PartRem[2][3] ),
	.A(n56), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U98 (
	.Y(n48),
	.A(a[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U99 (
	.Y(n29),
	.B(quotient[7]),
	.A(n49), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U100 (
	.Y(n30),
	.B(n29),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR2XLM U101 (
	.Y(n49),
	.B(a[7]),
	.A(\u_div/BInv [0]), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U102 (
	.Y(n54),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][4] ),
	.A(n44), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U103 (
	.Y(n56),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][2] ),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2XLM U104 (
	.Y(n55),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][3] ),
	.A(n42), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2XLM U105 (
	.Y(\u_div/PartRem[1][6] ),
	.S0(quotient[1]),
	.B(n60),
	.A(n54), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U106 (
	.Y(n60),
	.A(\u_div/SumTmp[1][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2XLM U107 (
	.Y(\u_div/PartRem[1][4] ),
	.S0(quotient[1]),
	.B(n69),
	.A(n56), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U108 (
	.Y(n69),
	.A(\u_div/SumTmp[1][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U109 (
	.Y(n39),
	.S0(quotient[4]),
	.B(\u_div/SumTmp[4][3] ),
	.A(n43), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U110 (
	.Y(\u_div/PartRem[2][6] ),
	.A(n53), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U111 (
	.Y(\u_div/PartRem[2][5] ),
	.A(n54), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2XLM U112 (
	.Y(\u_div/PartRem[1][7] ),
	.S0(quotient[1]),
	.B(n59),
	.A(n53), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U113 (
	.Y(n59),
	.A(\u_div/SumTmp[1][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U114 (
	.Y(n44),
	.S0(quotient[3]),
	.B(\u_div/SumTmp[3][3] ),
	.A(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2XLM U115 (
	.Y(n45),
	.S0(quotient[3]),
	.B(\u_div/SumTmp[3][4] ),
	.A(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2XLM U116 (
	.Y(n77),
	.B(\u_div/BInv [5]),
	.A(n91), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U117 (
	.Y(n64),
	.A(a[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U118 (
	.Y(n46),
	.B(\u_div/BInv [2]),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2XLM U119 (
	.Y(\u_div/PartRem[1][5] ),
	.S0(quotient[1]),
	.B(n63),
	.A(n55), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U120 (
	.Y(n63),
	.A(\u_div/SumTmp[1][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U121 (
	.Y(n75),
	.A(\u_div/SumTmp[1][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U122 (
	.Y(\u_div/PartRem[2][4] ),
	.A(n55), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U123 (
	.Y(\u_div/CryTmp[0][1] ),
	.B(FE_PT1_n92),
	.A(b[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U125 (
	.Y(\u_div/BInv [5]),
	.A(b[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR2XLM U127 (
	.Y(n50),
	.B(a[1]),
	.A(\u_div/BInv [0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U128 (
	.Y(\u_div/BInv [4]),
	.A(b[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U129 (
	.Y(\u_div/BInv [6]),
	.A(b[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U130 (
	.Y(n53),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][5] ),
	.A(n45), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X3M U131 (
	.Y(\u_div/PartRem[1][2] ),
	.S0(quotient[1]),
	.B(n79),
	.A(n58), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U132 (
	.Y(n71),
	.A(\u_div/SumTmp[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_2_0  (
	.S(\u_div/SumTmp[2][0] ),
	.CO(\u_div/CryTmp[2][1] ),
	.CI(HTIE_LTIEHI_NET),
	.B(\u_div/BInv [0]),
	.A(a[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_3_0  (
	.S(\u_div/SumTmp[3][0] ),
	.CO(\u_div/CryTmp[3][1] ),
	.CI(HTIE_LTIEHI_NET),
	.B(\u_div/BInv [0]),
	.A(a[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_4_0  (
	.S(\u_div/SumTmp[4][0] ),
	.CO(\u_div/CryTmp[4][1] ),
	.CI(HTIE_LTIEHI_NET),
	.B(\u_div/BInv [0]),
	.A(a[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_5_0  (
	.S(\u_div/SumTmp[5][0] ),
	.CO(\u_div/CryTmp[5][1] ),
	.CI(HTIE_LTIEHI_NET),
	.B(\u_div/BInv [0]),
	.A(a[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_6_0  (
	.S(\u_div/SumTmp[6][0] ),
	.CO(\u_div/CryTmp[6][1] ),
	.CI(HTIE_LTIEHI_NET),
	.B(\u_div/BInv [0]),
	.A(a[6]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SYS_CTRL_test_1 (
	RX_D_VLD, 
	RX_P_Data, 
	ALU_OUT, 
	OUT_Valid, 
	RdData, 
	RdData_Valid, 
	CLK, 
	RST, 
	fifo_full, 
	busyFall, 
	ALU_EN, 
	ALU_FUNC, 
	CLK_EN, 
	Address, 
	WrEn, 
	RdEn, 
	WrData, 
	TX_P_Data, 
	TX_D_VLD, 
	clk_div_en, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN1_rst_from_sync1, 
	VDD, 
	VSS);
   input RX_D_VLD;
   input [7:0] RX_P_Data;
   input [15:0] ALU_OUT;
   input OUT_Valid;
   input [7:0] RdData;
   input RdData_Valid;
   input CLK;
   input RST;
   input fifo_full;
   input busyFall;
   output ALU_EN;
   output [3:0] ALU_FUNC;
   output CLK_EN;
   output [3:0] Address;
   output WrEn;
   output RdEn;
   output [7:0] WrData;
   output [7:0] TX_P_Data;
   output TX_D_VLD;
   output clk_div_en;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN1_rst_from_sync1;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN13_SI_3_;
   wire FE_PHN12_SI_3_;
   wire LTIE_LTIELO_NET;
   wire FE_OFN4_reg_address_3_;
   wire FE_OFN3_reg_address_2_;
   wire N164;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n54;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire [3:0] current_state;
   wire [3:0] next_state;
   wire [3:0] address_;

   assign test_so = current_state[3] ;

   // Module instantiations
   DLY4X1M FE_PHC13_SI_3_ (
	.Y(FE_PHN13_SI_3_),
	.A(FE_PHN12_SI_3_), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC12_SI_3_ (
	.Y(FE_PHN12_SI_3_),
	.A(test_si), 
	.VDD(VDD), 
	.VSS(VSS));
   TIELOM LTIE_LTIELO (
	.Y(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M FE_OFC4_reg_address_3_ (
	.Y(Address[3]),
	.A(FE_OFN4_reg_address_3_), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M FE_OFC3_reg_address_2_ (
	.Y(Address[2]),
	.A(FE_OFN3_reg_address_2_), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \address__reg[3]  (
	.SI(address_[2]),
	.SE(test_se),
	.RN(RST),
	.Q(address_[3]),
	.D(n74),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \address__reg[2]  (
	.SI(address_[1]),
	.SE(test_se),
	.RN(RST),
	.Q(address_[2]),
	.D(n75),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \address__reg[1]  (
	.SI(address_[0]),
	.SE(test_se),
	.RN(RST),
	.Q(address_[1]),
	.D(n76),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \address__reg[0]  (
	.SI(FE_PHN13_SI_3_),
	.SE(test_se),
	.RN(FE_OFN1_rst_from_sync1),
	.Q(address_[0]),
	.D(n77),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[1]  (
	.SI(current_state[0]),
	.SE(test_se),
	.RN(FE_OFN1_rst_from_sync1),
	.Q(current_state[1]),
	.D(next_state[1]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[3]  (
	.SI(current_state[2]),
	.SE(test_se),
	.RN(FE_OFN1_rst_from_sync1),
	.Q(current_state[3]),
	.D(next_state[3]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[2]  (
	.SI(current_state[1]),
	.SE(test_se),
	.RN(FE_OFN1_rst_from_sync1),
	.Q(current_state[2]),
	.D(next_state[2]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[0]  (
	.SI(address_[3]),
	.SE(test_se),
	.RN(FE_OFN1_rst_from_sync1),
	.Q(current_state[0]),
	.D(next_state[0]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U13 (
	.Y(FE_OFN4_reg_address_3_),
	.B1(n26),
	.B0(n56),
	.A1N(address_[3]),
	.A0(n50), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U14 (
	.Y(n57),
	.B(n50),
	.A(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U15 (
	.Y(FE_OFN3_reg_address_2_),
	.B1(n25),
	.B0(n56),
	.A1N(address_[2]),
	.A0(n50), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U16 (
	.Y(n33),
	.B(n79),
	.A(n81), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U17 (
	.Y(n56),
	.B(RdEn),
	.A(n42), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X2M U18 (
	.Y(n42),
	.C(n83),
	.B(n80),
	.A(n41), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U19 (
	.Y(WrData[0]),
	.B(n22),
	.A(n57), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U20 (
	.Y(WrData[1]),
	.B(n24),
	.A(n57), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U21 (
	.Y(WrData[2]),
	.B(n25),
	.A(n57), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U22 (
	.Y(WrData[3]),
	.B(n26),
	.A(n57), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U23 (
	.Y(WrData[4]),
	.B(n27),
	.A(n57), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U24 (
	.Y(WrData[5]),
	.B(n28),
	.A(n57), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U25 (
	.Y(WrData[6]),
	.B(n54),
	.A(n57), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U26 (
	.Y(WrData[7]),
	.B(n78),
	.A(n57), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U27 (
	.Y(n35),
	.B(n55),
	.A(n53), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U28 (
	.Y(TX_D_VLD),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U29 (
	.Y(next_state[2]),
	.C(n34),
	.B(n33),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U30 (
	.Y(n34),
	.C0(n36),
	.B1(n35),
	.B0(n23),
	.A1(n20),
	.A0(RdEn), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U31 (
	.Y(n23),
	.A(n38), 
	.VDD(VDD), 
	.VSS(VSS));
   AND4X2M U32 (
	.Y(n36),
	.D(n35),
	.C(n37),
	.B(n22),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U33 (
	.Y(n81),
	.A(n51), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U34 (
	.Y(n79),
	.A(n70), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U35 (
	.Y(n43),
	.C(n52),
	.B(n27),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U36 (
	.Y(n82),
	.A(n55), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U37 (
	.Y(ALU_FUNC[2]),
	.B(n25),
	.A(n71), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U38 (
	.Y(ALU_FUNC[0]),
	.B(n22),
	.A(n71), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U39 (
	.Y(ALU_FUNC[3]),
	.B(n26),
	.A(n71), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U40 (
	.Y(ALU_FUNC[1]),
	.B(n24),
	.A(n71), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U41 (
	.Y(ALU_EN),
	.A(n68), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U42 (
	.Y(CLK_EN),
	.B(n30),
	.A(n68), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U43 (
	.Y(Address[0]),
	.C0(n70),
	.B1(n84),
	.B0(n50),
	.A1(n22),
	.A0(n56), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U44 (
	.Y(n84),
	.A(address_[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U45 (
	.Y(n41),
	.B(current_state[3]),
	.AN(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X2M U46 (
	.Y(RdEn),
	.C(n80),
	.B(current_state[2]),
	.A(n73), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U47 (
	.Y(n50),
	.C(current_state[0]),
	.B(n83),
	.A(n41), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U48 (
	.Y(n73),
	.B(current_state[1]),
	.A(current_state[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U49 (
	.Y(n83),
	.A(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U50 (
	.Y(n80),
	.A(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U51 (
	.Y(n69),
	.C(current_state[0]),
	.B(current_state[2]),
	.A(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U52 (
	.Y(Address[1]),
	.B1(n24),
	.B0(n56),
	.A1N(address_[1]),
	.A0(n50), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U53 (
	.Y(n55),
	.C(n73),
	.B(n83),
	.A(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U54 (
	.Y(n30),
	.B(n69),
	.A(current_state[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U55 (
	.Y(TX_P_Data[1]),
	.B1(n30),
	.B0(n66),
	.A1(n24),
	.A0(n55), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U56 (
	.Y(n66),
	.C1(n60),
	.C0(ALU_OUT[1]),
	.B1(n59),
	.B0(ALU_OUT[9]),
	.A1(RdData_Valid),
	.A0(RdData[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U57 (
	.Y(TX_P_Data[2]),
	.B1(n30),
	.B0(n65),
	.A1(n25),
	.A0(n55), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U58 (
	.Y(n65),
	.C1(n60),
	.C0(ALU_OUT[2]),
	.B1(n59),
	.B0(ALU_OUT[10]),
	.A1(RdData_Valid),
	.A0(RdData[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U59 (
	.Y(TX_P_Data[3]),
	.B1(n30),
	.B0(n64),
	.A1(n55),
	.A0(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U60 (
	.Y(n64),
	.C1(n60),
	.C0(ALU_OUT[3]),
	.B1(n59),
	.B0(ALU_OUT[11]),
	.A1(RdData_Valid),
	.A0(RdData[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U61 (
	.Y(TX_P_Data[4]),
	.B1(n30),
	.B0(n63),
	.A1(n27),
	.A0(n55), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U62 (
	.Y(n63),
	.C1(n60),
	.C0(ALU_OUT[4]),
	.B1(n59),
	.B0(ALU_OUT[12]),
	.A1(RdData_Valid),
	.A0(RdData[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U63 (
	.Y(TX_P_Data[5]),
	.B1(n30),
	.B0(n62),
	.A1(n28),
	.A0(n55), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U64 (
	.Y(n62),
	.C1(n60),
	.C0(ALU_OUT[5]),
	.B1(n59),
	.B0(ALU_OUT[13]),
	.A1(RdData_Valid),
	.A0(RdData[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U65 (
	.Y(TX_P_Data[6]),
	.B1(n30),
	.B0(n61),
	.A1(n54),
	.A0(n55), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U66 (
	.Y(n61),
	.C1(n60),
	.C0(ALU_OUT[6]),
	.B1(n59),
	.B0(ALU_OUT[14]),
	.A1(RdData_Valid),
	.A0(RdData[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U67 (
	.Y(TX_P_Data[7]),
	.B1(n30),
	.B0(n58),
	.A1(n55),
	.A0(n78), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U68 (
	.Y(n58),
	.C1(n60),
	.C0(ALU_OUT[7]),
	.B1(n59),
	.B0(ALU_OUT[15]),
	.A1(RdData[7]),
	.A0(RdData_Valid), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U69 (
	.Y(n60),
	.B(RdData_Valid),
	.AN(OUT_Valid), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U70 (
	.Y(n59),
	.B(RdData_Valid),
	.A(OUT_Valid), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U71 (
	.Y(n51),
	.C(n73),
	.B(current_state[0]),
	.A(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U72 (
	.Y(n25),
	.A(RX_P_Data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U73 (
	.Y(n24),
	.A(RX_P_Data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U74 (
	.Y(n70),
	.C(current_state[2]),
	.B(n80),
	.A(n41), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U75 (
	.Y(n22),
	.A(RX_P_Data[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U76 (
	.Y(n26),
	.A(RX_P_Data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U77 (
	.Y(WrEn),
	.B0(n33),
	.A1(n50),
	.A0(N164), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U78 (
	.Y(n74),
	.B0(Address[3]),
	.A1(n56),
	.A0(address_[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U79 (
	.Y(n77),
	.B1(address_[0]),
	.B0(n56),
	.A1N(n56),
	.A0(Address[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U80 (
	.Y(n75),
	.B0(Address[2]),
	.A1(address_[2]),
	.A0(n56), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U81 (
	.Y(n52),
	.D(RX_P_Data[6]),
	.C(RX_P_Data[2]),
	.B(n24),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U82 (
	.Y(n37),
	.D(RX_P_Data[5]),
	.C(RX_P_Data[1]),
	.B(n25),
	.A(n54), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI31X1M U83 (
	.Y(next_state[3]),
	.B0(n31),
	.A2(n30),
	.A1(RdData_Valid),
	.A0(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U84 (
	.Y(n31),
	.B0(RX_D_VLD),
	.A1(RdEn),
	.A0(ALU_EN), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U85 (
	.Y(n48),
	.C(current_state[2]),
	.B(current_state[3]),
	.A(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U86 (
	.Y(n68),
	.C(current_state[2]),
	.B(n41),
	.A(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U87 (
	.Y(n32),
	.B0(n11),
	.A1(ALU_EN),
	.A0(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   AND4X2M U88 (
	.Y(n11),
	.D(n37),
	.C(n35),
	.B(RX_P_Data[0]),
	.A(RX_P_Data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U89 (
	.Y(n49),
	.B0(RX_D_VLD),
	.A1(n51),
	.A0(n50), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U90 (
	.Y(n53),
	.B(RX_P_Data[3]),
	.A(RX_P_Data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U91 (
	.Y(n38),
	.C(n52),
	.B(RX_P_Data[0]),
	.A(RX_P_Data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2BB1X2M U92 (
	.Y(n47),
	.B0(n30),
	.A1N(RdData_Valid),
	.A0N(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U93 (
	.Y(next_state[0]),
	.D(n46),
	.C(n45),
	.B(n44),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U94 (
	.Y(n44),
	.B(n53),
	.A(n82), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U95 (
	.Y(n45),
	.B0(n49),
	.A2(n35),
	.A1(n38),
	.A0(n43), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI31X1M U96 (
	.Y(n46),
	.B0(RX_D_VLD),
	.A2(n48),
	.A1(n79),
	.A0(n47), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U97 (
	.Y(n28),
	.A(RX_P_Data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U98 (
	.Y(n54),
	.A(RX_P_Data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U99 (
	.Y(n27),
	.A(RX_P_Data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U100 (
	.Y(next_state[1]),
	.C(n40),
	.B(n32),
	.A(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U101 (
	.Y(n39),
	.B1(RX_D_VLD),
	.B0(n81),
	.A1(n35),
	.A0(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X2M U102 (
	.Y(n40),
	.C0(n42),
	.B0(n79),
	.A1(n20),
	.A0(n41), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U103 (
	.Y(n21),
	.A(n43), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U104 (
	.Y(n78),
	.A(RX_P_Data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U105 (
	.Y(n29),
	.B(OUT_Valid),
	.AN(fifo_full), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U106 (
	.Y(n20),
	.A(RX_D_VLD), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U107 (
	.Y(n76),
	.B0(Address[1]),
	.A1(address_[1]),
	.A0(n56), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X2M U108 (
	.Y(n71),
	.C(n72),
	.B(n56),
	.A(n57), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U109 (
	.Y(n72),
	.C(n69),
	.B(current_state[3]),
	.A(n82), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U110 (
	.Y(n67),
	.C1(n60),
	.C0(ALU_OUT[0]),
	.B1(n59),
	.B0(ALU_OUT[8]),
	.A1(RdData_Valid),
	.A0(RdData[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U111 (
	.Y(TX_P_Data[0]),
	.B1(n30),
	.B0(n67),
	.A1(n22),
	.A0(n55), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U112 (
	.Y(n12),
	.B(address_[0]),
	.AN(RX_P_Data[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U113 (
	.Y(n19),
	.B1(n12),
	.B0(RX_P_Data[1]),
	.A1N(address_[1]),
	.A0(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U114 (
	.Y(n13),
	.B(RX_P_Data[0]),
	.AN(address_[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U115 (
	.Y(n18),
	.B1(n13),
	.B0(address_[1]),
	.A1N(RX_P_Data[1]),
	.A0(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U116 (
	.Y(n15),
	.B(address_[2]),
	.A(RX_P_Data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U117 (
	.Y(n14),
	.B(address_[3]),
	.A(RX_P_Data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U118 (
	.Y(n17),
	.B(n14),
	.A(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U119 (
	.Y(n16),
	.D(RX_P_Data[4]),
	.C(RX_P_Data[5]),
	.B(RX_P_Data[6]),
	.A(RX_P_Data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND4X1M U120 (
	.Y(N164),
	.D(n16),
	.C(n17),
	.B(n18),
	.A(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U3 (
	.Y(clk_div_en),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module FIFO_test_1 (
	W_CLK, 
	W_RST, 
	W_INC, 
	R_CLK, 
	R_RST, 
	R_INC, 
	WR_DATA, 
	RD_DATA, 
	full, 
	empty, 
	test_si2, 
	test_si1, 
	test_so2, 
	test_so1, 
	test_se, 
	tx_clock__L3_N1, 
	tx_clock__L3_N2, 
	ref_clock__L5_N2, 
	ref_clock__L5_N3, 
	VDD, 
	VSS);
   input W_CLK;
   input W_RST;
   input W_INC;
   input R_CLK;
   input R_RST;
   input R_INC;
   input [7:0] WR_DATA;
   output [7:0] RD_DATA;
   output full;
   output empty;
   input test_si2;
   input test_si1;
   output test_so2;
   output test_so1;
   input test_se;
   input tx_clock__L3_N1;
   input tx_clock__L3_N2;
   input ref_clock__L5_N2;
   input ref_clock__L5_N3;
   inout VDD;
   inout VSS;

   // Internal wires
   wire empty_tx_valid;
   wire n1;
   wire [2:0] write_address;
   wire [2:0] read_address;
   wire [3:0] read_ptr_synch;
   wire [3:0] write_ptr;
   wire [3:0] read_ptr;
   wire [3:0] write_ptr_synch;

   assign test_so2 = write_ptr_synch[3] ;
   assign test_so1 = write_ptr_synch[0] ;

   // Module instantiations
   INVX2M U1 (
	.Y(empty),
	.A(empty_tx_valid), 
	.VDD(VDD), 
	.VSS(VSS));
   Ram_test_1 mem (
	.write_data({ WR_DATA[7],
		WR_DATA[6],
		WR_DATA[5],
		WR_DATA[4],
		WR_DATA[3],
		WR_DATA[2],
		WR_DATA[1],
		WR_DATA[0] }),
	.w_inc(W_INC),
	.r_inc(R_INC),
	.full(full),
	.empty(empty_tx_valid),
	.wraddress({ write_address[2],
		write_address[1],
		write_address[0] }),
	.rdaddress({ read_address[2],
		read_address[1],
		read_address[0] }),
	.clk(W_CLK),
	.rclk(R_CLK),
	.read_data({ RD_DATA[7],
		RD_DATA[6],
		RD_DATA[5],
		RD_DATA[4],
		RD_DATA[3],
		RD_DATA[2],
		RD_DATA[1],
		RD_DATA[0] }),
	.test_so(n1),
	.test_se(test_se),
	.ref_clock__L5_N2(ref_clock__L5_N2),
	.ref_clock__L5_N3(ref_clock__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   FIFO_Full_test_1 fifo_w (
	.wclk(W_CLK),
	.w_inc(W_INC),
	.r_inc(R_INC),
	.wrst_n(W_RST),
	.synch_readptr({ read_ptr_synch[3],
		read_ptr_synch[2],
		read_ptr_synch[1],
		read_ptr_synch[0] }),
	.full(full),
	.wraddress({ write_address[2],
		write_address[1],
		write_address[0] }),
	.write_ptr({ write_ptr[3],
		write_ptr[2],
		write_ptr[1],
		write_ptr[0] }),
	.test_si(empty_tx_valid),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   Synchronizer_test_0 read_synch (
	.pointer({ read_ptr[3],
		read_ptr[2],
		read_ptr[1],
		read_ptr[0] }),
	.clk(W_CLK),
	.rst(W_RST),
	.synchronized_pointer({ read_ptr_synch[3],
		read_ptr_synch[2],
		read_ptr_synch[1],
		read_ptr_synch[0] }),
	.test_si(n1),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   FIFO_Empty_test_1 fifo_rd (
	.rclk(tx_clock__L3_N1),
	.r_inc(R_INC),
	.w_inc(W_INC),
	.rrst_n(R_RST),
	.synch_wptr({ write_ptr_synch[3],
		write_ptr_synch[2],
		write_ptr_synch[1],
		write_ptr_synch[0] }),
	.empty(empty_tx_valid),
	.raddress({ read_address[2],
		read_address[1],
		read_address[0] }),
	.read_ptr({ read_ptr[3],
		read_ptr[2],
		read_ptr[1],
		read_ptr[0] }),
	.test_si(test_si1),
	.test_se(test_se),
	.tx_clock__L3_N2(tx_clock__L3_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   Synchronizer_test_1 write_synch (
	.pointer({ write_ptr[3],
		write_ptr[2],
		write_ptr[1],
		write_ptr[0] }),
	.clk(R_CLK),
	.rst(R_RST),
	.synchronized_pointer({ write_ptr_synch[3],
		write_ptr_synch[2],
		write_ptr_synch[1],
		write_ptr_synch[0] }),
	.test_si2(test_si2),
	.test_si1(read_ptr_synch[3]),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module Ram_test_1 (
	write_data, 
	w_inc, 
	r_inc, 
	full, 
	empty, 
	wraddress, 
	rdaddress, 
	clk, 
	rclk, 
	read_data, 
	test_so, 
	test_se, 
	ref_clock__L5_N2, 
	ref_clock__L5_N3, 
	VDD, 
	VSS);
   input [7:0] write_data;
   input w_inc;
   input r_inc;
   input full;
   input empty;
   input [2:0] wraddress;
   input [2:0] rdaddress;
   input clk;
   input rclk;
   output [7:0] read_data;
   output test_so;
   input test_se;
   input ref_clock__L5_N2;
   input ref_clock__L5_N3;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N9;
   wire N10;
   wire N11;
   wire \mem[0][7] ;
   wire \mem[0][6] ;
   wire \mem[0][5] ;
   wire \mem[0][4] ;
   wire \mem[0][3] ;
   wire \mem[0][2] ;
   wire \mem[0][1] ;
   wire \mem[0][0] ;
   wire \mem[1][7] ;
   wire \mem[1][6] ;
   wire \mem[1][5] ;
   wire \mem[1][4] ;
   wire \mem[1][3] ;
   wire \mem[1][2] ;
   wire \mem[1][1] ;
   wire \mem[1][0] ;
   wire \mem[2][7] ;
   wire \mem[2][6] ;
   wire \mem[2][5] ;
   wire \mem[2][4] ;
   wire \mem[2][3] ;
   wire \mem[2][2] ;
   wire \mem[2][1] ;
   wire \mem[2][0] ;
   wire \mem[3][7] ;
   wire \mem[3][6] ;
   wire \mem[3][5] ;
   wire \mem[3][4] ;
   wire \mem[3][3] ;
   wire \mem[3][2] ;
   wire \mem[3][1] ;
   wire \mem[3][0] ;
   wire \mem[4][7] ;
   wire \mem[4][6] ;
   wire \mem[4][5] ;
   wire \mem[4][4] ;
   wire \mem[4][3] ;
   wire \mem[4][2] ;
   wire \mem[4][1] ;
   wire \mem[4][0] ;
   wire \mem[5][7] ;
   wire \mem[5][6] ;
   wire \mem[5][5] ;
   wire \mem[5][4] ;
   wire \mem[5][3] ;
   wire \mem[5][2] ;
   wire \mem[5][1] ;
   wire \mem[5][0] ;
   wire \mem[6][7] ;
   wire \mem[6][6] ;
   wire \mem[6][5] ;
   wire \mem[6][4] ;
   wire \mem[6][3] ;
   wire \mem[6][2] ;
   wire \mem[6][1] ;
   wire \mem[6][0] ;
   wire \mem[7][7] ;
   wire \mem[7][6] ;
   wire \mem[7][5] ;
   wire \mem[7][4] ;
   wire \mem[7][3] ;
   wire \mem[7][2] ;
   wire \mem[7][1] ;
   wire \mem[7][0] ;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;
   wire n102;
   wire n103;
   wire n104;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n116;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;
   wire n165;
   wire n166;
   wire n167;
   wire n168;
   wire n169;
   wire n170;
   wire n171;
   wire n172;
   wire n173;
   wire n174;
   wire n176;
   wire n177;
   wire n178;

   assign N9 = rdaddress[0] ;
   assign N10 = rdaddress[1] ;
   assign N11 = rdaddress[2] ;
   assign test_so = \mem[7][7]  ;

   // Module instantiations
   SDFFQX2M \mem_reg[1][7]  (
	.SI(\mem[1][6] ),
	.SE(n176),
	.Q(\mem[1][7] ),
	.D(n141),
	.CK(ref_clock__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[1][6]  (
	.SI(\mem[1][5] ),
	.SE(n178),
	.Q(\mem[1][6] ),
	.D(n140),
	.CK(ref_clock__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[1][5]  (
	.SI(\mem[1][4] ),
	.SE(n177),
	.Q(\mem[1][5] ),
	.D(n139),
	.CK(ref_clock__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[1][4]  (
	.SI(\mem[1][3] ),
	.SE(n176),
	.Q(\mem[1][4] ),
	.D(n138),
	.CK(ref_clock__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[1][3]  (
	.SI(\mem[1][2] ),
	.SE(n178),
	.Q(\mem[1][3] ),
	.D(n137),
	.CK(ref_clock__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[1][2]  (
	.SI(\mem[1][1] ),
	.SE(n177),
	.Q(\mem[1][2] ),
	.D(n136),
	.CK(ref_clock__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[1][1]  (
	.SI(\mem[1][0] ),
	.SE(n176),
	.Q(\mem[1][1] ),
	.D(n135),
	.CK(ref_clock__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[1][0]  (
	.SI(\mem[0][7] ),
	.SE(n178),
	.Q(\mem[1][0] ),
	.D(n134),
	.CK(ref_clock__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[5][6]  (
	.SI(\mem[5][5] ),
	.SE(n177),
	.Q(\mem[5][6] ),
	.D(n108),
	.CK(ref_clock__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[5][5]  (
	.SI(\mem[5][4] ),
	.SE(n176),
	.Q(\mem[5][5] ),
	.D(n107),
	.CK(ref_clock__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[5][4]  (
	.SI(\mem[5][3] ),
	.SE(n178),
	.Q(\mem[5][4] ),
	.D(n106),
	.CK(ref_clock__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[5][3]  (
	.SI(\mem[5][2] ),
	.SE(n177),
	.Q(\mem[5][3] ),
	.D(n105),
	.CK(ref_clock__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[5][2]  (
	.SI(\mem[5][1] ),
	.SE(n176),
	.Q(\mem[5][2] ),
	.D(n104),
	.CK(ref_clock__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[5][1]  (
	.SI(\mem[5][0] ),
	.SE(n178),
	.Q(\mem[5][1] ),
	.D(n103),
	.CK(ref_clock__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[5][0]  (
	.SI(\mem[4][7] ),
	.SE(n177),
	.Q(\mem[5][0] ),
	.D(n102),
	.CK(ref_clock__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[3][7]  (
	.SI(\mem[3][6] ),
	.SE(n176),
	.Q(\mem[3][7] ),
	.D(n125),
	.CK(ref_clock__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[3][6]  (
	.SI(\mem[3][5] ),
	.SE(n178),
	.Q(\mem[3][6] ),
	.D(n124),
	.CK(ref_clock__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[3][5]  (
	.SI(\mem[3][4] ),
	.SE(n177),
	.Q(\mem[3][5] ),
	.D(n123),
	.CK(ref_clock__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[3][4]  (
	.SI(\mem[3][3] ),
	.SE(n176),
	.Q(\mem[3][4] ),
	.D(n122),
	.CK(ref_clock__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[3][3]  (
	.SI(\mem[3][2] ),
	.SE(n178),
	.Q(\mem[3][3] ),
	.D(n121),
	.CK(ref_clock__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[3][2]  (
	.SI(\mem[3][1] ),
	.SE(n177),
	.Q(\mem[3][2] ),
	.D(n120),
	.CK(ref_clock__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[3][1]  (
	.SI(\mem[3][0] ),
	.SE(n176),
	.Q(\mem[3][1] ),
	.D(n119),
	.CK(ref_clock__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[3][0]  (
	.SI(\mem[2][7] ),
	.SE(n178),
	.Q(\mem[3][0] ),
	.D(n118),
	.CK(ref_clock__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[7][7]  (
	.SI(\mem[7][6] ),
	.SE(n177),
	.Q(\mem[7][7] ),
	.D(n93),
	.CK(ref_clock__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[7][6]  (
	.SI(\mem[7][5] ),
	.SE(n176),
	.Q(\mem[7][6] ),
	.D(n92),
	.CK(ref_clock__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[7][5]  (
	.SI(\mem[7][4] ),
	.SE(n178),
	.Q(\mem[7][5] ),
	.D(n91),
	.CK(ref_clock__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[7][4]  (
	.SI(\mem[7][3] ),
	.SE(n177),
	.Q(\mem[7][4] ),
	.D(n90),
	.CK(ref_clock__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[7][3]  (
	.SI(\mem[7][2] ),
	.SE(n176),
	.Q(\mem[7][3] ),
	.D(n89),
	.CK(ref_clock__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[7][2]  (
	.SI(\mem[7][1] ),
	.SE(n178),
	.Q(\mem[7][2] ),
	.D(n88),
	.CK(ref_clock__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[7][1]  (
	.SI(\mem[7][0] ),
	.SE(n177),
	.Q(\mem[7][1] ),
	.D(n87),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[7][0]  (
	.SI(\mem[6][7] ),
	.SE(n176),
	.Q(\mem[7][0] ),
	.D(n86),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[2][7]  (
	.SI(\mem[2][6] ),
	.SE(n178),
	.Q(\mem[2][7] ),
	.D(n133),
	.CK(ref_clock__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[2][6]  (
	.SI(\mem[2][5] ),
	.SE(n177),
	.Q(\mem[2][6] ),
	.D(n132),
	.CK(ref_clock__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[2][5]  (
	.SI(\mem[2][4] ),
	.SE(n176),
	.Q(\mem[2][5] ),
	.D(n131),
	.CK(ref_clock__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[2][4]  (
	.SI(\mem[2][3] ),
	.SE(n178),
	.Q(\mem[2][4] ),
	.D(n130),
	.CK(ref_clock__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[2][3]  (
	.SI(\mem[2][2] ),
	.SE(n177),
	.Q(\mem[2][3] ),
	.D(n129),
	.CK(ref_clock__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[2][2]  (
	.SI(\mem[2][1] ),
	.SE(n176),
	.Q(\mem[2][2] ),
	.D(n128),
	.CK(ref_clock__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[2][1]  (
	.SI(\mem[2][0] ),
	.SE(n178),
	.Q(\mem[2][1] ),
	.D(n127),
	.CK(ref_clock__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[2][0]  (
	.SI(\mem[1][7] ),
	.SE(n177),
	.Q(\mem[2][0] ),
	.D(n126),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[6][7]  (
	.SI(\mem[6][6] ),
	.SE(n176),
	.Q(\mem[6][7] ),
	.D(n101),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[6][6]  (
	.SI(\mem[6][5] ),
	.SE(n178),
	.Q(\mem[6][6] ),
	.D(n100),
	.CK(ref_clock__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[6][5]  (
	.SI(\mem[6][4] ),
	.SE(n177),
	.Q(\mem[6][5] ),
	.D(n99),
	.CK(ref_clock__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[6][4]  (
	.SI(\mem[6][3] ),
	.SE(n176),
	.Q(\mem[6][4] ),
	.D(n98),
	.CK(ref_clock__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[6][3]  (
	.SI(\mem[6][2] ),
	.SE(n178),
	.Q(\mem[6][3] ),
	.D(n97),
	.CK(ref_clock__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[6][2]  (
	.SI(\mem[6][1] ),
	.SE(n177),
	.Q(\mem[6][2] ),
	.D(n96),
	.CK(ref_clock__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[6][1]  (
	.SI(\mem[6][0] ),
	.SE(n176),
	.Q(\mem[6][1] ),
	.D(n95),
	.CK(ref_clock__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[6][0]  (
	.SI(\mem[5][7] ),
	.SE(n178),
	.Q(\mem[6][0] ),
	.D(n94),
	.CK(ref_clock__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[0][7]  (
	.SI(\mem[0][6] ),
	.SE(n177),
	.Q(\mem[0][7] ),
	.D(n149),
	.CK(ref_clock__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[0][6]  (
	.SI(\mem[0][5] ),
	.SE(n176),
	.Q(\mem[0][6] ),
	.D(n148),
	.CK(ref_clock__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[0][5]  (
	.SI(\mem[0][4] ),
	.SE(n178),
	.Q(\mem[0][5] ),
	.D(n147),
	.CK(ref_clock__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[0][4]  (
	.SI(\mem[0][3] ),
	.SE(n177),
	.Q(\mem[0][4] ),
	.D(n146),
	.CK(ref_clock__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[0][3]  (
	.SI(\mem[0][2] ),
	.SE(n176),
	.Q(\mem[0][3] ),
	.D(n145),
	.CK(ref_clock__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[0][2]  (
	.SI(\mem[0][1] ),
	.SE(n178),
	.Q(\mem[0][2] ),
	.D(n144),
	.CK(ref_clock__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[0][1]  (
	.SI(\mem[0][0] ),
	.SE(n177),
	.Q(\mem[0][1] ),
	.D(n143),
	.CK(ref_clock__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[0][0]  (
	.SI(full),
	.SE(n176),
	.Q(\mem[0][0] ),
	.D(n142),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[4][7]  (
	.SI(\mem[4][6] ),
	.SE(n178),
	.Q(\mem[4][7] ),
	.D(n117),
	.CK(ref_clock__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[4][6]  (
	.SI(\mem[4][5] ),
	.SE(n177),
	.Q(\mem[4][6] ),
	.D(n116),
	.CK(ref_clock__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[4][5]  (
	.SI(\mem[4][4] ),
	.SE(n176),
	.Q(\mem[4][5] ),
	.D(n115),
	.CK(ref_clock__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[4][4]  (
	.SI(\mem[4][3] ),
	.SE(n178),
	.Q(\mem[4][4] ),
	.D(n114),
	.CK(ref_clock__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[4][3]  (
	.SI(\mem[4][2] ),
	.SE(n177),
	.Q(\mem[4][3] ),
	.D(n113),
	.CK(ref_clock__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[4][2]  (
	.SI(\mem[4][1] ),
	.SE(n176),
	.Q(\mem[4][2] ),
	.D(n112),
	.CK(ref_clock__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[4][1]  (
	.SI(\mem[4][0] ),
	.SE(n178),
	.Q(\mem[4][1] ),
	.D(n111),
	.CK(ref_clock__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX2M \mem_reg[4][0]  (
	.SI(\mem[3][7] ),
	.SE(n177),
	.Q(\mem[4][0] ),
	.D(n110),
	.CK(ref_clock__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFQX1M \mem_reg[5][7]  (
	.SI(\mem[5][6] ),
	.SE(n176),
	.Q(\mem[5][7] ),
	.D(n109),
	.CK(ref_clock__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U72 (
	.Y(n79),
	.C(n76),
	.B(n166),
	.A(n165), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U73 (
	.Y(n85),
	.C(n82),
	.B(n166),
	.A(n165), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U74 (
	.Y(n82),
	.B(wraddress[2]),
	.AN(n80), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U75 (
	.Y(n168),
	.A(write_data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U76 (
	.Y(n169),
	.A(write_data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U77 (
	.Y(n170),
	.A(write_data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U78 (
	.Y(n171),
	.A(write_data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U79 (
	.Y(n172),
	.A(write_data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U80 (
	.Y(n173),
	.A(write_data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U81 (
	.Y(n174),
	.A(write_data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U82 (
	.Y(n167),
	.A(write_data[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U83 (
	.Y(n142),
	.B1(n85),
	.B0(n167),
	.A1N(n85),
	.A0N(\mem[0][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U84 (
	.Y(n143),
	.B1(n85),
	.B0(n168),
	.A1N(n85),
	.A0N(\mem[0][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U85 (
	.Y(n144),
	.B1(n85),
	.B0(n169),
	.A1N(n85),
	.A0N(\mem[0][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U86 (
	.Y(n145),
	.B1(n85),
	.B0(n170),
	.A1N(n85),
	.A0N(\mem[0][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U87 (
	.Y(n146),
	.B1(n85),
	.B0(n171),
	.A1N(n85),
	.A0N(\mem[0][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U88 (
	.Y(n147),
	.B1(n85),
	.B0(n172),
	.A1N(n85),
	.A0N(\mem[0][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U89 (
	.Y(n148),
	.B1(n85),
	.B0(n173),
	.A1N(n85),
	.A0N(\mem[0][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U90 (
	.Y(n149),
	.B1(n85),
	.B0(n174),
	.A1N(n85),
	.A0N(\mem[0][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U91 (
	.Y(n110),
	.B1(n79),
	.B0(n167),
	.A1N(n79),
	.A0N(\mem[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U92 (
	.Y(n111),
	.B1(n79),
	.B0(n168),
	.A1N(n79),
	.A0N(\mem[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U93 (
	.Y(n112),
	.B1(n79),
	.B0(n169),
	.A1N(n79),
	.A0N(\mem[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U94 (
	.Y(n113),
	.B1(n79),
	.B0(n170),
	.A1N(n79),
	.A0N(\mem[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U95 (
	.Y(n114),
	.B1(n79),
	.B0(n171),
	.A1N(n79),
	.A0N(\mem[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U96 (
	.Y(n115),
	.B1(n79),
	.B0(n172),
	.A1N(n79),
	.A0N(\mem[4][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U97 (
	.Y(n116),
	.B1(n79),
	.B0(n173),
	.A1N(n79),
	.A0N(\mem[4][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U98 (
	.Y(n117),
	.B1(n79),
	.B0(n174),
	.A1N(n79),
	.A0N(\mem[4][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U99 (
	.Y(n94),
	.B1(n77),
	.B0(n167),
	.A1N(n77),
	.A0N(\mem[6][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U100 (
	.Y(n102),
	.B1(n78),
	.B0(n167),
	.A1N(n78),
	.A0N(\mem[5][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U101 (
	.Y(n118),
	.B1(n81),
	.B0(n167),
	.A1N(n81),
	.A0N(\mem[3][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U102 (
	.Y(n126),
	.B1(n83),
	.B0(n167),
	.A1N(n83),
	.A0N(\mem[2][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U103 (
	.Y(n134),
	.B1(n84),
	.B0(n167),
	.A1N(n84),
	.A0N(\mem[1][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U104 (
	.Y(n86),
	.B1(n167),
	.B0(n75),
	.A1N(n75),
	.A0N(\mem[7][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U106 (
	.Y(n75),
	.C(wraddress[1]),
	.B(n76),
	.A(wraddress[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U107 (
	.Y(n87),
	.B1(n168),
	.B0(n75),
	.A1N(n75),
	.A0N(\mem[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U108 (
	.Y(n88),
	.B1(n169),
	.B0(n75),
	.A1N(n75),
	.A0N(\mem[7][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U109 (
	.Y(n89),
	.B1(n170),
	.B0(n75),
	.A1N(n75),
	.A0N(\mem[7][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U110 (
	.Y(n90),
	.B1(n171),
	.B0(n75),
	.A1N(n75),
	.A0N(\mem[7][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U111 (
	.Y(n91),
	.B1(n172),
	.B0(n75),
	.A1N(n75),
	.A0N(\mem[7][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U112 (
	.Y(n92),
	.B1(n173),
	.B0(n75),
	.A1N(n75),
	.A0N(\mem[7][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U113 (
	.Y(n93),
	.B1(n174),
	.B0(n75),
	.A1N(n75),
	.A0N(\mem[7][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U114 (
	.Y(n95),
	.B1(n77),
	.B0(n168),
	.A1N(n77),
	.A0N(\mem[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U115 (
	.Y(n96),
	.B1(n77),
	.B0(n169),
	.A1N(n77),
	.A0N(\mem[6][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U116 (
	.Y(n97),
	.B1(n77),
	.B0(n170),
	.A1N(n77),
	.A0N(\mem[6][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U117 (
	.Y(n98),
	.B1(n77),
	.B0(n171),
	.A1N(n77),
	.A0N(\mem[6][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U118 (
	.Y(n99),
	.B1(n77),
	.B0(n172),
	.A1N(n77),
	.A0N(\mem[6][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U119 (
	.Y(n100),
	.B1(n77),
	.B0(n173),
	.A1N(n77),
	.A0N(\mem[6][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U120 (
	.Y(n101),
	.B1(n77),
	.B0(n174),
	.A1N(n77),
	.A0N(\mem[6][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U121 (
	.Y(n103),
	.B1(n78),
	.B0(n168),
	.A1N(n78),
	.A0N(\mem[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U122 (
	.Y(n104),
	.B1(n78),
	.B0(n169),
	.A1N(n78),
	.A0N(\mem[5][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U123 (
	.Y(n105),
	.B1(n78),
	.B0(n170),
	.A1N(n78),
	.A0N(\mem[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U124 (
	.Y(n106),
	.B1(n78),
	.B0(n171),
	.A1N(n78),
	.A0N(\mem[5][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U125 (
	.Y(n107),
	.B1(n78),
	.B0(n172),
	.A1N(n78),
	.A0N(\mem[5][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U126 (
	.Y(n108),
	.B1(n78),
	.B0(n173),
	.A1N(n78),
	.A0N(\mem[5][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U127 (
	.Y(n109),
	.B1(n78),
	.B0(n174),
	.A1N(n78),
	.A0N(\mem[5][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U128 (
	.Y(n119),
	.B1(n81),
	.B0(n168),
	.A1N(n81),
	.A0N(\mem[3][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U129 (
	.Y(n120),
	.B1(n81),
	.B0(n169),
	.A1N(n81),
	.A0N(\mem[3][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U130 (
	.Y(n121),
	.B1(n81),
	.B0(n170),
	.A1N(n81),
	.A0N(\mem[3][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U131 (
	.Y(n122),
	.B1(n81),
	.B0(n171),
	.A1N(n81),
	.A0N(\mem[3][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U132 (
	.Y(n123),
	.B1(n81),
	.B0(n172),
	.A1N(n81),
	.A0N(\mem[3][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U133 (
	.Y(n124),
	.B1(n81),
	.B0(n173),
	.A1N(n81),
	.A0N(\mem[3][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U134 (
	.Y(n125),
	.B1(n81),
	.B0(n174),
	.A1N(n81),
	.A0N(\mem[3][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U135 (
	.Y(n127),
	.B1(n83),
	.B0(n168),
	.A1N(n83),
	.A0N(\mem[2][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U136 (
	.Y(n128),
	.B1(n83),
	.B0(n169),
	.A1N(n83),
	.A0N(\mem[2][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U137 (
	.Y(n129),
	.B1(n83),
	.B0(n170),
	.A1N(n83),
	.A0N(\mem[2][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U138 (
	.Y(n130),
	.B1(n83),
	.B0(n171),
	.A1N(n83),
	.A0N(\mem[2][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U139 (
	.Y(n131),
	.B1(n83),
	.B0(n172),
	.A1N(n83),
	.A0N(\mem[2][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U140 (
	.Y(n132),
	.B1(n83),
	.B0(n173),
	.A1N(n83),
	.A0N(\mem[2][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U141 (
	.Y(n133),
	.B1(n83),
	.B0(n174),
	.A1N(n83),
	.A0N(\mem[2][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U142 (
	.Y(n135),
	.B1(n84),
	.B0(n168),
	.A1N(n84),
	.A0N(\mem[1][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U143 (
	.Y(n136),
	.B1(n84),
	.B0(n169),
	.A1N(n84),
	.A0N(\mem[1][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U144 (
	.Y(n137),
	.B1(n84),
	.B0(n170),
	.A1N(n84),
	.A0N(\mem[1][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U145 (
	.Y(n138),
	.B1(n84),
	.B0(n171),
	.A1N(n84),
	.A0N(\mem[1][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U146 (
	.Y(n139),
	.B1(n84),
	.B0(n172),
	.A1N(n84),
	.A0N(\mem[1][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U147 (
	.Y(n140),
	.B1(n84),
	.B0(n173),
	.A1N(n84),
	.A0N(\mem[1][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U148 (
	.Y(n141),
	.B1(n84),
	.B0(n174),
	.A1N(n84),
	.A0N(\mem[1][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U149 (
	.Y(n80),
	.B(full),
	.AN(w_inc), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U150 (
	.Y(n76),
	.B(n80),
	.A(wraddress[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U151 (
	.Y(n78),
	.C(wraddress[0]),
	.B(n166),
	.A(n76), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U152 (
	.Y(n77),
	.C(wraddress[1]),
	.B(n165),
	.A(n76), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U153 (
	.Y(n81),
	.C(n82),
	.B(wraddress[0]),
	.A(wraddress[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U154 (
	.Y(n84),
	.C(n82),
	.B(n166),
	.A(wraddress[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U155 (
	.Y(n83),
	.C(n82),
	.B(n165),
	.A(wraddress[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U156 (
	.Y(n165),
	.A(wraddress[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U157 (
	.Y(n166),
	.A(wraddress[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U158 (
	.Y(read_data[0]),
	.S0(N11),
	.B(n66),
	.A(n67), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U159 (
	.Y(n67),
	.S1(N10),
	.S0(n158),
	.D(\mem[3][0] ),
	.C(\mem[2][0] ),
	.B(\mem[1][0] ),
	.A(\mem[0][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U160 (
	.Y(n66),
	.S1(N10),
	.S0(n157),
	.D(\mem[7][0] ),
	.C(\mem[6][0] ),
	.B(\mem[5][0] ),
	.A(\mem[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U161 (
	.Y(read_data[1]),
	.S0(N11),
	.B(n68),
	.A(n69), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U162 (
	.Y(n69),
	.S1(N10),
	.S0(n158),
	.D(\mem[3][1] ),
	.C(\mem[2][1] ),
	.B(\mem[1][1] ),
	.A(\mem[0][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U163 (
	.Y(n68),
	.S1(N10),
	.S0(n157),
	.D(\mem[7][1] ),
	.C(\mem[6][1] ),
	.B(\mem[5][1] ),
	.A(\mem[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U164 (
	.Y(read_data[2]),
	.S0(N11),
	.B(n70),
	.A(n71), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U165 (
	.Y(n71),
	.S1(N10),
	.S0(n158),
	.D(\mem[3][2] ),
	.C(\mem[2][2] ),
	.B(\mem[1][2] ),
	.A(\mem[0][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U166 (
	.Y(n70),
	.S1(N10),
	.S0(n157),
	.D(\mem[7][2] ),
	.C(\mem[6][2] ),
	.B(\mem[5][2] ),
	.A(\mem[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U167 (
	.Y(read_data[3]),
	.S0(N11),
	.B(n72),
	.A(n73), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U168 (
	.Y(n73),
	.S1(N10),
	.S0(n158),
	.D(\mem[3][3] ),
	.C(\mem[2][3] ),
	.B(\mem[1][3] ),
	.A(\mem[0][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U169 (
	.Y(n72),
	.S1(N10),
	.S0(n157),
	.D(\mem[7][3] ),
	.C(\mem[6][3] ),
	.B(\mem[5][3] ),
	.A(\mem[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U170 (
	.Y(read_data[4]),
	.S0(N11),
	.B(n74),
	.A(n150), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U171 (
	.Y(n150),
	.S1(N10),
	.S0(n158),
	.D(\mem[3][4] ),
	.C(\mem[2][4] ),
	.B(\mem[1][4] ),
	.A(\mem[0][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U172 (
	.Y(n74),
	.S1(N10),
	.S0(n157),
	.D(\mem[7][4] ),
	.C(\mem[6][4] ),
	.B(\mem[5][4] ),
	.A(\mem[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U173 (
	.Y(read_data[5]),
	.S0(N11),
	.B(n151),
	.A(n152), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U174 (
	.Y(n152),
	.S1(N10),
	.S0(n158),
	.D(\mem[3][5] ),
	.C(\mem[2][5] ),
	.B(\mem[1][5] ),
	.A(\mem[0][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U175 (
	.Y(n151),
	.S1(N10),
	.S0(n157),
	.D(\mem[7][5] ),
	.C(\mem[6][5] ),
	.B(\mem[5][5] ),
	.A(\mem[4][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U176 (
	.Y(read_data[6]),
	.S0(N11),
	.B(n153),
	.A(n154), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U177 (
	.Y(n154),
	.S1(N10),
	.S0(n158),
	.D(\mem[3][6] ),
	.C(\mem[2][6] ),
	.B(\mem[1][6] ),
	.A(\mem[0][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U178 (
	.Y(n153),
	.S1(N10),
	.S0(n157),
	.D(\mem[7][6] ),
	.C(\mem[6][6] ),
	.B(\mem[5][6] ),
	.A(\mem[4][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U179 (
	.Y(read_data[7]),
	.S0(N11),
	.B(n155),
	.A(n156), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U180 (
	.Y(n156),
	.S1(N10),
	.S0(n158),
	.D(\mem[3][7] ),
	.C(\mem[2][7] ),
	.B(\mem[1][7] ),
	.A(\mem[0][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U181 (
	.Y(n155),
	.S1(N10),
	.S0(n157),
	.D(\mem[7][7] ),
	.C(\mem[6][7] ),
	.B(\mem[5][7] ),
	.A(\mem[4][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U182 (
	.Y(n157),
	.A(N9), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U183 (
	.Y(n158),
	.A(N9), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X4M U184 (
	.Y(n176),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X4M U185 (
	.Y(n177),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X4M U186 (
	.Y(n178),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module FIFO_Full_test_1 (
	wclk, 
	w_inc, 
	r_inc, 
	wrst_n, 
	synch_readptr, 
	full, 
	wraddress, 
	write_ptr, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input wclk;
   input w_inc;
   input r_inc;
   input wrst_n;
   input [3:0] synch_readptr;
   output full;
   output [2:0] wraddress;
   output [3:0] write_ptr;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;

   // Module instantiations
   SDFFRQX2M full_reg (
	.SI(write_ptr[3]),
	.SE(test_se),
	.RN(wrst_n),
	.Q(full),
	.D(n20),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \bin_cnt_reg[3]  (
	.SI(wraddress[2]),
	.SE(test_se),
	.RN(wrst_n),
	.Q(write_ptr[3]),
	.D(n21),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \bin_cnt_reg[2]  (
	.SI(wraddress[1]),
	.SE(test_se),
	.RN(wrst_n),
	.Q(wraddress[2]),
	.D(n22),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \bin_cnt_reg[1]  (
	.SI(wraddress[0]),
	.SE(test_se),
	.RN(wrst_n),
	.Q(wraddress[1]),
	.D(n23),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U9 (
	.Y(n15),
	.B(n9),
	.A(w_inc), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U10 (
	.Y(n16),
	.B(synch_readptr[1]),
	.A(write_ptr[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U11 (
	.Y(write_ptr[0]),
	.B(wraddress[1]),
	.A(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U12 (
	.Y(n14),
	.B(n8),
	.A(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U13 (
	.Y(n22),
	.B(n13),
	.A(wraddress[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U14 (
	.Y(n21),
	.B(n12),
	.A(write_ptr[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U15 (
	.Y(n12),
	.B(wraddress[2]),
	.AN(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U16 (
	.Y(n9),
	.D(n19),
	.C(n18),
	.B(n17),
	.A(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U17 (
	.Y(n19),
	.B(synch_readptr[3]),
	.A(write_ptr[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U18 (
	.Y(n17),
	.B(synch_readptr[0]),
	.A(write_ptr[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U19 (
	.Y(n18),
	.B(write_ptr[2]),
	.A(synch_readptr[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U20 (
	.Y(n13),
	.B(wraddress[1]),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U21 (
	.Y(write_ptr[2]),
	.B(wraddress[2]),
	.A(write_ptr[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U22 (
	.Y(write_ptr[1]),
	.B(wraddress[2]),
	.A(wraddress[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U23 (
	.Y(n23),
	.B(n14),
	.A(wraddress[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI31X1M U24 (
	.Y(n20),
	.B0(n11),
	.A2(n10),
	.A1(r_inc),
	.A0(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U25 (
	.Y(n11),
	.B(n10),
	.A(full), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U26 (
	.Y(n10),
	.B(r_inc),
	.A(w_inc), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U27 (
	.Y(n24),
	.B(n15),
	.A(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \bin_cnt_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(wrst_n),
	.QN(n8),
	.Q(wraddress[0]),
	.D(n24),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module Synchronizer_test_0 (
	pointer, 
	clk, 
	rst, 
	synchronized_pointer, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input [3:0] pointer;
   input clk;
   input rst;
   output [3:0] synchronized_pointer;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire [3:0] internal_pointer;

   // Module instantiations
   SDFFRQX2M \synchronized_pointer_reg[1]  (
	.SI(synchronized_pointer[0]),
	.SE(test_se),
	.RN(rst),
	.Q(synchronized_pointer[1]),
	.D(internal_pointer[1]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \synchronized_pointer_reg[0]  (
	.SI(internal_pointer[3]),
	.SE(test_se),
	.RN(rst),
	.Q(synchronized_pointer[0]),
	.D(internal_pointer[0]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \synchronized_pointer_reg[3]  (
	.SI(synchronized_pointer[2]),
	.SE(test_se),
	.RN(rst),
	.Q(synchronized_pointer[3]),
	.D(internal_pointer[3]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \synchronized_pointer_reg[2]  (
	.SI(synchronized_pointer[1]),
	.SE(test_se),
	.RN(rst),
	.Q(synchronized_pointer[2]),
	.D(internal_pointer[2]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \internal_pointer_reg[3]  (
	.SI(internal_pointer[2]),
	.SE(test_se),
	.RN(rst),
	.Q(internal_pointer[3]),
	.D(pointer[3]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \internal_pointer_reg[2]  (
	.SI(internal_pointer[1]),
	.SE(test_se),
	.RN(rst),
	.Q(internal_pointer[2]),
	.D(pointer[2]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \internal_pointer_reg[1]  (
	.SI(internal_pointer[0]),
	.SE(test_se),
	.RN(rst),
	.Q(internal_pointer[1]),
	.D(pointer[1]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \internal_pointer_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(rst),
	.Q(internal_pointer[0]),
	.D(pointer[0]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module FIFO_Empty_test_1 (
	rclk, 
	r_inc, 
	w_inc, 
	rrst_n, 
	synch_wptr, 
	empty, 
	raddress, 
	read_ptr, 
	test_si, 
	test_se, 
	tx_clock__L3_N2, 
	VDD, 
	VSS);
   input rclk;
   input r_inc;
   input w_inc;
   input rrst_n;
   input [3:0] synch_wptr;
   output empty;
   output [2:0] raddress;
   output [3:0] read_ptr;
   input test_si;
   input test_se;
   input tx_clock__L3_N2;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N7;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n11;
   wire n13;
   wire n15;
   wire n17;
   wire n2;

   // Module instantiations
   SDFFRQX2M \bin_cnt_reg[3]  (
	.SI(raddress[2]),
	.SE(test_se),
	.RN(rrst_n),
	.Q(read_ptr[3]),
	.D(n11),
	.CK(rclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \bin_cnt_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(rrst_n),
	.Q(raddress[0]),
	.D(n17),
	.CK(tx_clock__L3_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \bin_cnt_reg[2]  (
	.SI(raddress[1]),
	.SE(test_se),
	.RN(rrst_n),
	.Q(raddress[2]),
	.D(n13),
	.CK(tx_clock__L3_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX4M \bin_cnt_reg[1]  (
	.SI(raddress[0]),
	.SE(test_se),
	.RN(rrst_n),
	.Q(raddress[1]),
	.D(n15),
	.CK(tx_clock__L3_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSQX1M empty_reg (
	.SN(rrst_n),
	.SI(read_ptr[3]),
	.SE(test_se),
	.Q(empty),
	.D(N7),
	.CK(rclk), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U4 (
	.Y(n3),
	.B(n4),
	.AN(raddress[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U5 (
	.Y(N7),
	.D(n9),
	.C(n8),
	.B(n7),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U6 (
	.Y(n7),
	.B(read_ptr[3]),
	.A(synch_wptr[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U7 (
	.Y(n6),
	.B(read_ptr[2]),
	.A(synch_wptr[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U8 (
	.Y(n9),
	.B(read_ptr[1]),
	.A(synch_wptr[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U9 (
	.Y(n17),
	.B(n5),
	.A(raddress[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U10 (
	.Y(n15),
	.B(n4),
	.A(raddress[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U11 (
	.Y(n4),
	.B(raddress[0]),
	.AN(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U12 (
	.Y(n8),
	.B(read_ptr[0]),
	.A(synch_wptr[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U13 (
	.Y(n5),
	.B(r_inc),
	.AN(empty), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U14 (
	.Y(read_ptr[1]),
	.B(raddress[2]),
	.A(raddress[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U15 (
	.Y(read_ptr[0]),
	.B(raddress[1]),
	.A(raddress[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U16 (
	.Y(read_ptr[2]),
	.B(raddress[2]),
	.A(read_ptr[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U17 (
	.Y(n13),
	.B(n3),
	.A(raddress[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U18 (
	.Y(n11),
	.B(n2),
	.A(read_ptr[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U19 (
	.Y(n2),
	.B(raddress[2]),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module Synchronizer_test_1 (
	pointer, 
	clk, 
	rst, 
	synchronized_pointer, 
	test_si2, 
	test_si1, 
	test_se, 
	VDD, 
	VSS);
   input [3:0] pointer;
   input clk;
   input rst;
   output [3:0] synchronized_pointer;
   input test_si2;
   input test_si1;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN7_SI_0_;
   wire FE_PHN6_SI_0_;
   wire [3:0] internal_pointer;

   // Module instantiations
   DLY4X1M FE_PHC7_SI_0_ (
	.Y(FE_PHN7_SI_0_),
	.A(FE_PHN6_SI_0_), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC6_SI_0_ (
	.Y(FE_PHN6_SI_0_),
	.A(test_si2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \synchronized_pointer_reg[3]  (
	.SI(synchronized_pointer[2]),
	.SE(test_se),
	.RN(rst),
	.Q(synchronized_pointer[3]),
	.D(internal_pointer[3]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \synchronized_pointer_reg[2]  (
	.SI(synchronized_pointer[1]),
	.SE(test_se),
	.RN(rst),
	.Q(synchronized_pointer[2]),
	.D(internal_pointer[2]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \synchronized_pointer_reg[1]  (
	.SI(FE_PHN7_SI_0_),
	.SE(test_se),
	.RN(rst),
	.Q(synchronized_pointer[1]),
	.D(internal_pointer[1]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \synchronized_pointer_reg[0]  (
	.SI(internal_pointer[3]),
	.SE(test_se),
	.RN(rst),
	.Q(synchronized_pointer[0]),
	.D(internal_pointer[0]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \internal_pointer_reg[3]  (
	.SI(internal_pointer[2]),
	.SE(test_se),
	.RN(rst),
	.Q(internal_pointer[3]),
	.D(pointer[3]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \internal_pointer_reg[2]  (
	.SI(internal_pointer[1]),
	.SE(test_se),
	.RN(rst),
	.Q(internal_pointer[2]),
	.D(pointer[2]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \internal_pointer_reg[1]  (
	.SI(internal_pointer[0]),
	.SE(test_se),
	.RN(rst),
	.Q(internal_pointer[1]),
	.D(pointer[1]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \internal_pointer_reg[0]  (
	.SI(test_si1),
	.SE(test_se),
	.RN(rst),
	.Q(internal_pointer[0]),
	.D(pointer[0]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module UART_RX_test_1 (
	RX_IN, 
	Prescale, 
	PAR_EN, 
	PAR_TYP, 
	CLK, 
	RST, 
	P_DATA, 
	data_valid, 
	par_err, 
	stp_err, 
	test_si, 
	test_so, 
	test_se, 
	rx_clock__L3_N1, 
	rx_clock__L3_N2, 
	rx_clock__L3_N3, 
	VDD, 
	VSS);
   input RX_IN;
   input [5:0] Prescale;
   input PAR_EN;
   input PAR_TYP;
   input CLK;
   input RST;
   output [7:0] P_DATA;
   output data_valid;
   output par_err;
   output stp_err;
   input test_si;
   output test_so;
   input test_se;
   input rx_clock__L3_N1;
   input rx_clock__L3_N2;
   input rx_clock__L3_N3;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PT0_;
   wire FE_UNCONNECTED_0;
   wire disable_bit_cnt;
   wire data_sample_enable;
   wire sampled_bit;
   wire strt_glitch;
   wire start_check_en;
   wire stop_check_en;
   wire parity_check_en;
   wire deserial_enable;
   wire dis_err;
   wire parity_bit;
   wire n4;
   wire n5;
   wire n6;
   wire [2:0] bit_cnt;
   wire [5:0] edge_cnt;

   // Module instantiations
   edge_bit_counter_prescalar_width6_bit_width_count3_test_1 EDGE_U0 (
	.clk(rx_clock__L3_N1),
	.rst(RST),
	.prescale({ Prescale[5],
		Prescale[4],
		Prescale[3],
		Prescale[2],
		Prescale[1],
		Prescale[0] }),
	.enable(data_sample_enable),
	.disable_bit_count(disable_bit_cnt),
	.bit_count({ bit_cnt[2],
		bit_cnt[1],
		bit_cnt[0] }),
	.edge_count({ edge_cnt[5],
		edge_cnt[4],
		edge_cnt[3],
		edge_cnt[2],
		edge_cnt[1],
		edge_cnt[0] }),
	.test_si(test_si),
	.test_so(n6),
	.test_se(test_se),
	.rx_clock__L3_N2(rx_clock__L3_N2),
	.rx_clock__L3_N3(rx_clock__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   data_sampling_prescalar_WIDTH6_scaler6_test_1 sampling (
	.clk(rx_clock__L3_N2),
	.rst(RST),
	.edge_count({ edge_cnt[5],
		edge_cnt[4],
		edge_cnt[3],
		edge_cnt[2],
		edge_cnt[1],
		edge_cnt[0] }),
	.data_sample_en(data_sample_enable),
	.prescalar({ Prescale[5],
		Prescale[4],
		Prescale[3],
		Prescale[2],
		Prescale[1],
		Prescale[0] }),
	.RX_IN(RX_IN),
	.sampled_bit(sampled_bit),
	.test_si(n4),
	.test_so(test_so),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   FSM_RX_bit_count_width3_edge_cnt_width6_prescale_width6_test_1 controller (
	.RX_IN(RX_IN),
	.clk(CLK),
	.rst(RST),
	.parity_enable(PAR_EN),
	.bit_cnt({ bit_cnt[2],
		bit_cnt[1],
		bit_cnt[0] }),
	.edge_cnt({ edge_cnt[5],
		edge_cnt[4],
		edge_cnt[3],
		edge_cnt[2],
		edge_cnt[1],
		edge_cnt[0] }),
	.parity_error(par_err),
	.start_glitch(strt_glitch),
	.stop_error(stp_err),
	.Prescalar({ Prescale[5],
		Prescale[4],
		Prescale[3],
		Prescale[2],
		Prescale[1],
		Prescale[0] }),
	.dat_samp_en(data_sample_enable),
	.enable(FE_PT0_),
	.strt_chk_en(start_check_en),
	.stp_chk_en(stop_check_en),
	.par_chk_en(parity_check_en),
	.data_valid(data_valid),
	.des_en(deserial_enable),
	.disable_bit_count(disable_bit_cnt),
	.disable_parity_err(dis_err),
	.test_si(n6),
	.test_so(n5),
	.test_se(test_se),
	.rx_clock__L3_N1(rx_clock__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   deserializer_edge_width6_scaler_width6_data_width8_test_1 deserial (
	.clk(CLK),
	.rst(RST),
	.parity_type(PAR_TYP),
	.edge_count({ edge_cnt[5],
		edge_cnt[4],
		edge_cnt[3],
		edge_cnt[2],
		edge_cnt[1],
		edge_cnt[0] }),
	.prescale({ Prescale[5],
		Prescale[4],
		Prescale[3],
		Prescale[2],
		Prescale[1],
		Prescale[0] }),
	.sampled_bit(sampled_bit),
	.des_en(deserial_enable),
	.P_data({ P_DATA[7],
		P_DATA[6],
		P_DATA[5],
		P_DATA[4],
		P_DATA[3],
		P_DATA[2],
		P_DATA[1],
		P_DATA[0] }),
	.parity(parity_bit),
	.test_si(n5),
	.test_se(test_se),
	.rx_clock__L3_N1(rx_clock__L3_N1),
	.rx_clock__L3_N2(rx_clock__L3_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   parity_chk_test_1 par_checker (
	.clk(rx_clock__L3_N2),
	.rst(RST),
	.parity_bit(parity_bit),
	.disable_err(dis_err),
	.par_chk_en(parity_check_en),
	.sampled_bit(sampled_bit),
	.par_err(par_err),
	.test_so(n4),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   strt_chk start_checker (
	.sampled_bit(sampled_bit),
	.strt_chk_en(start_check_en),
	.strt_err(strt_glitch), 
	.VDD(VDD), 
	.VSS(VSS));
   stp_chk stop_checker (
	.sampled_bit(sampled_bit),
	.stp_chk_en(stop_check_en),
	.stp_chk_err(stp_err), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module edge_bit_counter_prescalar_width6_bit_width_count3_test_1 (
	clk, 
	rst, 
	prescale, 
	enable, 
	disable_bit_count, 
	bit_count, 
	edge_count, 
	test_si, 
	test_so, 
	test_se, 
	rx_clock__L3_N2, 
	rx_clock__L3_N3, 
	VDD, 
	VSS);
   input clk;
   input rst;
   input [5:0] prescale;
   input enable;
   input disable_bit_count;
   output [2:0] bit_count;
   output [5:0] edge_count;
   input test_si;
   output test_so;
   input test_se;
   input rx_clock__L3_N2;
   input rx_clock__L3_N3;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N9;
   wire N13;
   wire N14;
   wire N15;
   wire N16;
   wire N18;
   wire N19;
   wire N20;
   wire N21;
   wire N22;
   wire N23;
   wire N26;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire \add_20/carry[5] ;
   wire \add_20/carry[4] ;
   wire \add_20/carry[3] ;
   wire \add_20/carry[2] ;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n58;
   wire n59;
   wire [5:0] prescale_reg;

   assign test_so = prescale_reg[5] ;

   // Module instantiations
   SDFFRQX2M \bit_count_reg[2]  (
	.SI(n51),
	.SE(n59),
	.RN(rst),
	.Q(bit_count[2]),
	.D(n47),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \bit_count_reg[1]  (
	.SI(bit_count[0]),
	.SE(n59),
	.RN(rst),
	.Q(bit_count[1]),
	.D(n48),
	.CK(rx_clock__L3_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \bit_count_reg[0]  (
	.SI(test_si),
	.SE(n59),
	.RN(rst),
	.Q(bit_count[0]),
	.D(n49),
	.CK(rx_clock__L3_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \prescale_reg_reg[5]  (
	.SI(prescale_reg[4]),
	.SE(n59),
	.RN(rst),
	.Q(prescale_reg[5]),
	.D(prescale[5]),
	.CK(rx_clock__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \prescale_reg_reg[0]  (
	.SI(edge_count[5]),
	.SE(n59),
	.RN(rst),
	.Q(prescale_reg[0]),
	.D(prescale[0]),
	.CK(rx_clock__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \prescale_reg_reg[1]  (
	.SI(prescale_reg[0]),
	.SE(n59),
	.RN(rst),
	.Q(prescale_reg[1]),
	.D(prescale[1]),
	.CK(rx_clock__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \prescale_reg_reg[4]  (
	.SI(prescale_reg[3]),
	.SE(n59),
	.RN(rst),
	.Q(prescale_reg[4]),
	.D(prescale[4]),
	.CK(rx_clock__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \prescale_reg_reg[3]  (
	.SI(prescale_reg[2]),
	.SE(n59),
	.RN(rst),
	.Q(prescale_reg[3]),
	.D(prescale[3]),
	.CK(rx_clock__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \prescale_reg_reg[2]  (
	.SI(prescale_reg[1]),
	.SE(n59),
	.RN(rst),
	.Q(prescale_reg[2]),
	.D(prescale[2]),
	.CK(rx_clock__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \edge_count_reg[0]  (
	.SI(n52),
	.SE(n59),
	.RN(rst),
	.Q(edge_count[0]),
	.D(N18),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \edge_count_reg[5]  (
	.SI(edge_count[4]),
	.SE(n59),
	.RN(rst),
	.Q(edge_count[5]),
	.D(N23),
	.CK(rx_clock__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \edge_count_reg[1]  (
	.SI(edge_count[0]),
	.SE(n59),
	.RN(rst),
	.Q(edge_count[1]),
	.D(N19),
	.CK(rx_clock__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \edge_count_reg[4]  (
	.SI(n50),
	.SE(n59),
	.RN(rst),
	.Q(edge_count[4]),
	.D(N22),
	.CK(rx_clock__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \edge_count_reg[2]  (
	.SI(edge_count[1]),
	.SE(n59),
	.RN(rst),
	.Q(edge_count[2]),
	.D(N20),
	.CK(rx_clock__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \edge_count_reg[3]  (
	.SI(n27),
	.SE(n59),
	.RN(rst),
	.Q(edge_count[3]),
	.D(N21),
	.CK(rx_clock__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U6 (
	.Y(n26),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX2M U19 (
	.Y(n31),
	.C(N9),
	.B(n33),
	.AN(disable_bit_count), 
	.VDD(VDD), 
	.VSS(VSS));
   OR3X2M U20 (
	.Y(n32),
	.C(n26),
	.B(disable_bit_count),
	.A(N26), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U21 (
	.Y(n34),
	.D(n36),
	.C(n35),
	.B(N9),
	.A(enable), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U22 (
	.Y(n35),
	.B(n37),
	.A(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U23 (
	.Y(n37),
	.B0(n39),
	.A1(n53),
	.A0(n38), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U24 (
	.Y(N22),
	.B(n34),
	.AN(N16), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U25 (
	.Y(N21),
	.B(n34),
	.AN(N15), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U26 (
	.Y(N20),
	.B(n34),
	.AN(N14), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U27 (
	.Y(N19),
	.B(n34),
	.AN(N13), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI32X1M U28 (
	.Y(n47),
	.B1(n52),
	.B0(n29),
	.A2(n28),
	.A1(bit_count[2]),
	.A0(n51), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U29 (
	.Y(n52),
	.A(bit_count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U30 (
	.Y(n29),
	.B0(n30),
	.A1(n51),
	.A0(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U31 (
	.Y(n51),
	.A(bit_count[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U32 (
	.Y(n49),
	.B1(n31),
	.B0(bit_count[0]),
	.A1N(bit_count[0]),
	.A0(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U33 (
	.Y(n30),
	.B0(n32),
	.A1(n31),
	.A0(bit_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U34 (
	.Y(n48),
	.B1(n28),
	.B0(bit_count[1]),
	.A1N(bit_count[1]),
	.A0N(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U35 (
	.Y(n28),
	.B(n26),
	.A(bit_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI33X2M U36 (
	.Y(n45),
	.B2(n50),
	.B1(n27),
	.B0(n41),
	.A2(edge_count[3]),
	.A1(prescale[4]),
	.A0(n46), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U37 (
	.Y(n50),
	.A(edge_count[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI33X2M U38 (
	.Y(n46),
	.B2(prescale[3]),
	.B1(n55),
	.B0(edge_count[2]),
	.A2(prescale[2]),
	.A1(n54),
	.A0(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U39 (
	.Y(n27),
	.A(edge_count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U40 (
	.Y(n39),
	.D(prescale[4]),
	.C(prescale[3]),
	.B(prescale[2]),
	.A(n53), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U41 (
	.Y(n38),
	.B0(n41),
	.A1(n40),
	.A0(prescale[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U42 (
	.Y(n40),
	.B(prescale[3]),
	.A(n55), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U43 (
	.Y(n36),
	.B(prescale[0]),
	.A(prescale[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U44 (
	.Y(n53),
	.A(prescale[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U45 (
	.Y(n55),
	.A(prescale[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U46 (
	.Y(n54),
	.A(prescale[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U47 (
	.Y(n41),
	.C(prescale[4]),
	.B(n54),
	.A(n55), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U48 (
	.Y(N23),
	.B(n34),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U49 (
	.Y(n1),
	.B(edge_count[5]),
	.A(\add_20/carry[5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U50 (
	.Y(N18),
	.B(n34),
	.A(edge_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND4X2M U51 (
	.Y(n33),
	.D(n36),
	.C(n42),
	.B(edge_count[0]),
	.A(edge_count[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U52 (
	.Y(n42),
	.B0(edge_count[5]),
	.A1(n44),
	.A0(n43), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U53 (
	.Y(n44),
	.D(n39),
	.C(edge_count[2]),
	.B(edge_count[3]),
	.A(edge_count[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX2M U54 (
	.Y(n43),
	.C(n45),
	.B(n53),
	.AN(edge_count[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U55 (
	.S(N15),
	.CO(\add_20/carry[4] ),
	.B(\add_20/carry[3] ),
	.A(edge_count[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U56 (
	.S(N14),
	.CO(\add_20/carry[3] ),
	.B(\add_20/carry[2] ),
	.A(edge_count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U57 (
	.S(N13),
	.CO(\add_20/carry[2] ),
	.B(edge_count[0]),
	.A(edge_count[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U58 (
	.S(N16),
	.CO(\add_20/carry[5] ),
	.B(\add_20/carry[4] ),
	.A(edge_count[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U59 (
	.Y(n2),
	.B(prescale_reg[0]),
	.AN(prescale[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U60 (
	.Y(n25),
	.B1(n2),
	.B0(prescale[1]),
	.A1N(prescale_reg[1]),
	.A0(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U61 (
	.Y(n3),
	.B(prescale[0]),
	.AN(prescale_reg[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U62 (
	.Y(n24),
	.B1(n3),
	.B0(prescale_reg[1]),
	.A1N(prescale[1]),
	.A0(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U63 (
	.Y(n23),
	.B(prescale[5]),
	.A(prescale_reg[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U64 (
	.Y(n21),
	.B(prescale[4]),
	.A(prescale_reg[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U65 (
	.Y(n20),
	.B(prescale[2]),
	.A(prescale_reg[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U66 (
	.Y(n4),
	.B(prescale[3]),
	.A(prescale_reg[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X1M U67 (
	.Y(n22),
	.C(n4),
	.B(n20),
	.A(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X1M U68 (
	.Y(N26),
	.D(n22),
	.C(n23),
	.B(n24),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U69 (
	.Y(N9),
	.A(N26), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U70 (
	.Y(n58),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U71 (
	.Y(n59),
	.A(n58), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module data_sampling_prescalar_WIDTH6_scaler6_test_1 (
	clk, 
	rst, 
	edge_count, 
	data_sample_en, 
	prescalar, 
	RX_IN, 
	sampled_bit, 
	test_si, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input clk;
   input rst;
   input [5:0] edge_count;
   input data_sample_en;
   input [5:0] prescalar;
   input RX_IN;
   output sampled_bit;
   input test_si;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire conseq_sampled_bit;
   wire N8;
   wire N9;
   wire N10;
   wire N11;
   wire N12;
   wire N15;
   wire N16;
   wire N17;
   wire N18;
   wire N19;
   wire N20;
   wire N21;
   wire N34;
   wire N35;
   wire N36;
   wire n23;
   wire \add_31/carry[4] ;
   wire \add_31/carry[3] ;
   wire \add_31/carry[2] ;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire [1:0] sampled_count;

   assign test_so = sampled_count[1] ;

   // Module instantiations
   SDFFRQX2M conseq_sampled_bit_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(rst),
	.Q(conseq_sampled_bit),
	.D(N36),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sampled_count_reg[1]  (
	.SI(sampled_count[0]),
	.SE(test_se),
	.RN(rst),
	.Q(sampled_count[1]),
	.D(N35),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sampled_count_reg[0]  (
	.SI(sampled_bit),
	.SE(test_se),
	.RN(rst),
	.Q(sampled_count[0]),
	.D(N34),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M sampled_bit_reg (
	.SI(conseq_sampled_bit),
	.SE(test_se),
	.RN(rst),
	.Q(sampled_bit),
	.D(n23),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U6 (
	.Y(n1),
	.B(prescalar[1]),
	.A(prescalar[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U7 (
	.S(N9),
	.CO(\add_31/carry[3] ),
	.B(\add_31/carry[2] ),
	.A(prescalar[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U8 (
	.S(N10),
	.CO(\add_31/carry[4] ),
	.B(\add_31/carry[3] ),
	.A(prescalar[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U9 (
	.S(N8),
	.CO(\add_31/carry[2] ),
	.B(prescalar[1]),
	.A(prescalar[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U10 (
	.S(N11),
	.CO(N12),
	.B(\add_31/carry[4] ),
	.A(prescalar[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U12 (
	.Y(N15),
	.A(prescalar[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U13 (
	.Y(N16),
	.B0(n1),
	.A1N(prescalar[2]),
	.A0N(prescalar[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U14 (
	.Y(n2),
	.B(prescalar[3]),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U15 (
	.Y(N17),
	.B0(n2),
	.A1N(prescalar[3]),
	.A0N(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U16 (
	.Y(N18),
	.B(n2),
	.A(prescalar[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X1M U17 (
	.Y(N20),
	.C(n2),
	.B(prescalar[5]),
	.A(prescalar[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U18 (
	.Y(n3),
	.B0(prescalar[5]),
	.A1(n2),
	.A0(prescalar[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U19 (
	.Y(N19),
	.B(n3),
	.AN(N20), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U20 (
	.Y(n4),
	.B(N15),
	.AN(edge_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U21 (
	.Y(n7),
	.B1(n4),
	.B0(edge_count[1]),
	.A1N(N16),
	.A0(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U22 (
	.Y(n5),
	.B(edge_count[0]),
	.AN(N15), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U23 (
	.Y(n6),
	.B1(n5),
	.B0(N16),
	.A1N(edge_count[1]),
	.A0(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BBX1M U24 (
	.Y(n11),
	.D(n6),
	.C(n7),
	.BN(edge_count[5]),
	.AN(N20), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U25 (
	.Y(n10),
	.B(edge_count[4]),
	.A(N19), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U26 (
	.Y(n9),
	.B(edge_count[2]),
	.A(N17), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U27 (
	.Y(n8),
	.B(edge_count[3]),
	.A(N18), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U28 (
	.Y(N21),
	.D(n8),
	.C(n9),
	.B(n10),
	.A(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U29 (
	.Y(n23),
	.S0(conseq_sampled_bit),
	.B(sampled_count[1]),
	.A(sampled_bit), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U30 (
	.Y(N35),
	.B(n13),
	.A(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U31 (
	.Y(n13),
	.B(sampled_count[1]),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U32 (
	.Y(n14),
	.B(RX_IN),
	.A(sampled_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U33 (
	.Y(N34),
	.B(n19),
	.A(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U34 (
	.Y(n19),
	.B(sampled_count[0]),
	.A(RX_IN), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X1M U35 (
	.Y(n12),
	.B0(N36),
	.A1(data_sample_en),
	.A0(N21), 
	.VDD(VDD), 
	.VSS(VSS));
   OA21X1M U36 (
	.Y(N36),
	.B0(data_sample_en),
	.A1(n21),
	.A0(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U37 (
	.Y(n21),
	.D(n26),
	.C(n25),
	.B(n24),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U38 (
	.Y(n26),
	.B(N8),
	.A(edge_count[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U39 (
	.Y(n25),
	.B(N10),
	.A(edge_count[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U40 (
	.Y(n24),
	.B(N9),
	.A(edge_count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X1M U41 (
	.Y(n22),
	.C(n29),
	.B(n28),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U42 (
	.Y(n29),
	.B(N12),
	.A(edge_count[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U43 (
	.Y(n28),
	.B(N15),
	.A(edge_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U44 (
	.Y(n27),
	.B(N11),
	.A(edge_count[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U45 (
	.Y(n20),
	.D(n32),
	.C(edge_count[5]),
	.B(n31),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U46 (
	.Y(n32),
	.B(edge_count[0]),
	.A(prescalar[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U47 (
	.Y(n31),
	.B(edge_count[4]),
	.A(prescalar[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X1M U48 (
	.Y(n30),
	.C(n35),
	.B(n34),
	.A(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U49 (
	.Y(n35),
	.B(prescalar[3]),
	.A(edge_count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U50 (
	.Y(n34),
	.B(prescalar[4]),
	.A(edge_count[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U51 (
	.Y(n33),
	.B(prescalar[2]),
	.A(edge_count[1]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module FSM_RX_bit_count_width3_edge_cnt_width6_prescale_width6_test_1 (
	RX_IN, 
	clk, 
	rst, 
	parity_enable, 
	bit_cnt, 
	edge_cnt, 
	parity_error, 
	start_glitch, 
	stop_error, 
	Prescalar, 
	dat_samp_en, 
	enable, 
	strt_chk_en, 
	stp_chk_en, 
	par_chk_en, 
	data_valid, 
	des_en, 
	disable_bit_count, 
	disable_parity_err, 
	test_si, 
	test_so, 
	test_se, 
	rx_clock__L3_N1, 
	VDD, 
	VSS);
   input RX_IN;
   input clk;
   input rst;
   input parity_enable;
   input [2:0] bit_cnt;
   input [5:0] edge_cnt;
   input parity_error;
   input start_glitch;
   input stop_error;
   input [5:0] Prescalar;
   output dat_samp_en;
   output enable;
   output strt_chk_en;
   output stp_chk_en;
   output par_chk_en;
   output data_valid;
   output des_en;
   output disable_bit_count;
   output disable_parity_err;
   input test_si;
   output test_so;
   input test_se;
   input rx_clock__L3_N1;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N171;
   wire N172;
   wire N173;
   wire N174;
   wire N175;
   wire N176;
   wire N177;
   wire n52;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire \r111/EQ ;
   wire \r111/B[0] ;
   wire \r111/B[1] ;
   wire \r111/B[2] ;
   wire \r111/B[3] ;
   wire \r111/B[5] ;
   wire \r111/B[9] ;
   wire \add_223/carry[4] ;
   wire \add_223/carry[3] ;
   wire n2;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n53;
   wire n54;
   wire [5:0] prescale_reg;
   wire [2:0] current_state;
   wire [2:0] next_state;

   assign test_so = prescale_reg[5] ;

   // Module instantiations
   SDFFRQX2M \current_state_reg[2]  (
	.SI(n51),
	.SE(test_se),
	.RN(rst),
	.Q(current_state[2]),
	.D(next_state[2]),
	.CK(rx_clock__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(rst),
	.Q(current_state[0]),
	.D(next_state[0]),
	.CK(rx_clock__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[1]  (
	.SI(current_state[0]),
	.SE(test_se),
	.RN(rst),
	.Q(current_state[1]),
	.D(next_state[1]),
	.CK(rx_clock__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \prescale_reg_reg[5]  (
	.SI(prescale_reg[4]),
	.SE(test_se),
	.RN(rst),
	.Q(prescale_reg[5]),
	.D(Prescalar[5]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \prescale_reg_reg[1]  (
	.SI(\r111/B[0] ),
	.SE(test_se),
	.RN(rst),
	.Q(N171),
	.D(Prescalar[1]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \prescale_reg_reg[4]  (
	.SI(prescale_reg[3]),
	.SE(test_se),
	.RN(rst),
	.Q(prescale_reg[4]),
	.D(Prescalar[4]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \prescale_reg_reg[3]  (
	.SI(N172),
	.SE(test_se),
	.RN(rst),
	.Q(prescale_reg[3]),
	.D(Prescalar[3]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \prescale_reg_reg[0]  (
	.SI(n54),
	.SE(test_se),
	.RN(rst),
	.Q(prescale_reg[0]),
	.D(Prescalar[0]),
	.CK(rx_clock__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \prescale_reg_reg[2]  (
	.SI(N171),
	.SE(test_se),
	.RN(rst),
	.Q(prescale_reg[2]),
	.D(Prescalar[2]),
	.CK(rx_clock__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U14 (
	.Y(next_state[2]),
	.C1(n56),
	.C0(\r111/EQ ),
	.B1(n48),
	.B0(n58),
	.A1(n36),
	.A0(n57), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U15 (
	.Y(n36),
	.A(\r111/EQ ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3XLM U16 (
	.Y(n58),
	.C(\r111/EQ ),
	.B(n53),
	.A(n60), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B11X2M U17 (
	.Y(next_state[1]),
	.C0(n47),
	.B0(n59),
	.A1N(n58),
	.A0(n48), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4XLM U18 (
	.Y(n59),
	.D(n49),
	.C(n51),
	.B(n55),
	.A(\r111/EQ ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U19 (
	.Y(n47),
	.A(n63), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI32XLM U20 (
	.Y(n63),
	.B1(n57),
	.B0(\r111/EQ ),
	.A2(n53),
	.A1(n48),
	.A0(n64), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2XLM U21 (
	.Y(n64),
	.B(n60),
	.A(\r111/EQ ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U22 (
	.Y(n24),
	.A(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U23 (
	.Y(n66),
	.B(n50),
	.A(n67), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U24 (
	.Y(n48),
	.A(des_en), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U25 (
	.Y(disable_bit_count),
	.B(n50),
	.A(n66), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U26 (
	.Y(n26),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U27 (
	.Y(n25),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21XLM U28 (
	.Y(n65),
	.B0(\r111/EQ ),
	.A1(n49),
	.A0(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4XLM U29 (
	.Y(data_valid),
	.D(n36),
	.C(n56),
	.B(parity_error),
	.A(stop_error), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21BX2M U30 (
	.Y(n2),
	.B0N(n7),
	.A1(prescale_reg[4]),
	.A0(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X2M U31 (
	.Y(next_state[0]),
	.C0(n47),
	.B0(n62),
	.A1(n61),
	.A0(RX_IN), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U32 (
	.Y(n62),
	.C(n26),
	.B(n65),
	.A(n55), 
	.VDD(VDD), 
	.VSS(VSS));
   OA21X2M U33 (
	.Y(n61),
	.B0(n66),
	.A1(n56),
	.A0(n36), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U34 (
	.Y(n4),
	.B(prescale_reg[0]),
	.A(N171), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21BXLM U35 (
	.Y(n69),
	.B0N(N177),
	.A1(n52),
	.A0(\r111/EQ ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U36 (
	.Y(n22),
	.A(edge_cnt[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U37 (
	.Y(n23),
	.A(edge_cnt[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U38 (
	.Y(n21),
	.A(edge_cnt[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U39 (
	.Y(stp_chk_en),
	.B(n56),
	.A(n52), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U40 (
	.Y(des_en),
	.C(n51),
	.B(current_state[2]),
	.A(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U41 (
	.Y(n67),
	.B(current_state[0]),
	.A(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U42 (
	.Y(n56),
	.B(n67),
	.A(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U43 (
	.Y(n51),
	.A(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U44 (
	.Y(n60),
	.C(bit_cnt[0]),
	.B(bit_cnt[1]),
	.A(bit_cnt[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U45 (
	.Y(disable_parity_err),
	.B1(n68),
	.B0(current_state[1]),
	.A1(n51),
	.A0(n50), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U46 (
	.Y(n49),
	.A(start_glitch), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3BX2M U47 (
	.Y(strt_chk_en),
	.C(current_state[1]),
	.B(n52),
	.AN(n55), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U48 (
	.Y(par_chk_en),
	.B(n57),
	.A(n52), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U49 (
	.Y(n57),
	.B(n55),
	.A(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U50 (
	.Y(n50),
	.A(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U51 (
	.Y(n68),
	.B(n50),
	.A(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U52 (
	.Y(n55),
	.B(n50),
	.A(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U53 (
	.Y(n53),
	.A(parity_enable), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U54 (
	.Y(N172),
	.A(prescale_reg[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U56 (
	.Y(dat_samp_en),
	.B0(n56),
	.A1(n67),
	.A0(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U57 (
	.Y(N176),
	.B(prescale_reg[5]),
	.A(\add_223/carry[4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U58 (
	.Y(N175),
	.B(\add_223/carry[4] ),
	.A(prescale_reg[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U59 (
	.Y(\add_223/carry[4] ),
	.B(prescale_reg[4]),
	.A(\add_223/carry[3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U60 (
	.Y(N174),
	.B(\add_223/carry[3] ),
	.A(prescale_reg[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U61 (
	.Y(\add_223/carry[3] ),
	.B(prescale_reg[3]),
	.A(prescale_reg[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U62 (
	.Y(N173),
	.B(prescale_reg[2]),
	.A(prescale_reg[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U63 (
	.Y(\r111/B[0] ),
	.A(prescale_reg[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U64 (
	.Y(\r111/B[1] ),
	.B0(n4),
	.A1N(N171),
	.A0N(prescale_reg[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U65 (
	.Y(n5),
	.B(prescale_reg[2]),
	.A(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U66 (
	.Y(\r111/B[2] ),
	.B0(n5),
	.A1N(prescale_reg[2]),
	.A0N(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U67 (
	.Y(n6),
	.B(prescale_reg[3]),
	.A(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U68 (
	.Y(\r111/B[3] ),
	.B0(n6),
	.A1N(prescale_reg[3]),
	.A0N(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U69 (
	.Y(n7),
	.B(prescale_reg[4]),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U70 (
	.Y(\r111/B[9] ),
	.B(prescale_reg[5]),
	.A(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U71 (
	.Y(\r111/B[5] ),
	.B0(\r111/B[9] ),
	.A1(prescale_reg[5]),
	.A0(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U72 (
	.Y(n14),
	.B(\r111/B[3] ),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U73 (
	.Y(n13),
	.B(n2),
	.A(edge_cnt[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U74 (
	.Y(n8),
	.B(\r111/B[0] ),
	.AN(edge_cnt[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U75 (
	.Y(n9),
	.B1(n8),
	.B0(edge_cnt[1]),
	.A1N(\r111/B[1] ),
	.A0(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX1M U76 (
	.Y(n20),
	.C(n9),
	.B(n13),
	.AN(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U77 (
	.Y(n19),
	.B(\r111/B[2] ),
	.A(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U78 (
	.Y(n11),
	.B(\r111/B[0] ),
	.AN(edge_cnt[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2BB1X1M U79 (
	.Y(n10),
	.B0(\r111/B[1] ),
	.A1N(edge_cnt[1]),
	.A0N(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X1M U80 (
	.Y(n12),
	.C0(n10),
	.B0(n19),
	.A1(n11),
	.A0(edge_cnt[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U81 (
	.Y(n15),
	.C0(n12),
	.B1(n23),
	.B0(\r111/B[2] ),
	.A1(n22),
	.A0(\r111/B[3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI32X1M U82 (
	.Y(n16),
	.B1(n2),
	.B0(edge_cnt[4]),
	.A2(n24),
	.A1(n14),
	.A0(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U83 (
	.Y(n18),
	.B(\r111/B[5] ),
	.A(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U84 (
	.Y(n17),
	.C0(\r111/B[9] ),
	.B1(n21),
	.B0(\r111/B[5] ),
	.A1(n25),
	.A0(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U85 (
	.Y(\r111/EQ ),
	.D(n18),
	.C(n26),
	.B(n19),
	.A(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U86 (
	.Y(n27),
	.B(N171),
	.AN(edge_cnt[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U87 (
	.Y(n31),
	.B1(n27),
	.B0(edge_cnt[1]),
	.A1N(N172),
	.A0(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U88 (
	.Y(n28),
	.B(edge_cnt[0]),
	.AN(N171), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U89 (
	.Y(n30),
	.B1(n28),
	.B0(N172),
	.A1N(edge_cnt[1]),
	.A0(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U90 (
	.Y(n29),
	.B(edge_cnt[5]),
	.A(N176), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X1M U91 (
	.Y(n35),
	.C(n29),
	.B(n30),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U92 (
	.Y(n34),
	.B(edge_cnt[4]),
	.A(N175), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U93 (
	.Y(n33),
	.B(edge_cnt[2]),
	.A(N173), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U94 (
	.Y(n32),
	.B(edge_cnt[3]),
	.A(N174), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U95 (
	.Y(N177),
	.D(n32),
	.C(n33),
	.B(n34),
	.A(n35), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M flag_reg (
	.SI(n50),
	.SE(test_se),
	.RN(rst),
	.QN(n52),
	.Q(n54),
	.D(n69),
	.CK(rx_clock__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module deserializer_edge_width6_scaler_width6_data_width8_test_1 (
	clk, 
	rst, 
	parity_type, 
	edge_count, 
	prescale, 
	sampled_bit, 
	des_en, 
	P_data, 
	parity, 
	test_si, 
	test_se, 
	rx_clock__L3_N1, 
	rx_clock__L3_N2, 
	VDD, 
	VSS);
   input clk;
   input rst;
   input parity_type;
   input [5:0] edge_count;
   input [5:0] prescale;
   input sampled_bit;
   input des_en;
   output [7:0] P_data;
   output parity;
   input test_si;
   input test_se;
   input rx_clock__L3_N1;
   input rx_clock__L3_N2;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N3;
   wire N4;
   wire N5;
   wire N6;
   wire N7;
   wire N8;
   wire N9;
   wire N14;
   wire n5;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n20;
   wire n22;
   wire n24;
   wire n26;
   wire n28;
   wire n30;
   wire n32;
   wire n34;
   wire \add_17/carry[4] ;
   wire \add_17/carry[3] ;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;

   assign N3 = prescale[1] ;

   // Module instantiations
   SDFFRQX2M parity_reg (
	.SI(n12),
	.SE(test_se),
	.RN(rst),
	.Q(parity),
	.D(N14),
	.CK(rx_clock__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_data_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(rst),
	.Q(P_data[0]),
	.D(n20),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_data_reg[7]  (
	.SI(n13),
	.SE(test_se),
	.RN(rst),
	.Q(P_data[7]),
	.D(n34),
	.CK(rx_clock__L3_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_data_reg[5]  (
	.SI(n36),
	.SE(test_se),
	.RN(rst),
	.Q(P_data[5]),
	.D(n30),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_data_reg[4]  (
	.SI(n37),
	.SE(test_se),
	.RN(rst),
	.Q(P_data[4]),
	.D(n28),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_data_reg[3]  (
	.SI(n38),
	.SE(test_se),
	.RN(rst),
	.Q(P_data[3]),
	.D(n26),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_data_reg[1]  (
	.SI(P_data[0]),
	.SE(test_se),
	.RN(rst),
	.Q(P_data[1]),
	.D(n22),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_data_reg[6]  (
	.SI(n35),
	.SE(test_se),
	.RN(rst),
	.Q(P_data[6]),
	.D(n32),
	.CK(rx_clock__L3_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_data_reg[2]  (
	.SI(n39),
	.SE(test_se),
	.RN(rst),
	.Q(P_data[2]),
	.D(n24),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U3 (
	.Y(n22),
	.B1(n38),
	.B0(n5),
	.A1(n39),
	.A0(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U4 (
	.Y(n24),
	.B1(n37),
	.B0(n5),
	.A1(n38),
	.A0(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U5 (
	.Y(n26),
	.B1(n36),
	.B0(n5),
	.A1(n37),
	.A0(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U6 (
	.Y(n28),
	.B1(n35),
	.B0(n5),
	.A1(n36),
	.A0(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U7 (
	.Y(n30),
	.B1(n13),
	.B0(n5),
	.A1(n35),
	.A0(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U8 (
	.Y(n32),
	.B1(n12),
	.B0(n5),
	.A1(n13),
	.A0(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U9 (
	.Y(n11),
	.A(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U10 (
	.Y(n5),
	.B(N9),
	.A(des_en), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U11 (
	.Y(n20),
	.B1(n39),
	.B0(n5),
	.A1N(P_data[0]),
	.A0N(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U12 (
	.Y(n34),
	.B1(n12),
	.B0(n11),
	.A1N(n11),
	.A0N(sampled_bit), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U13 (
	.Y(N4),
	.A(prescale[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U14 (
	.Y(n17),
	.B(P_data[6]),
	.A(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U15 (
	.Y(N14),
	.C(parity_type),
	.B(n15),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U16 (
	.Y(n15),
	.C(n16),
	.B(P_data[0]),
	.A(P_data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U17 (
	.Y(n14),
	.C(n17),
	.B(n36),
	.A(n35), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U18 (
	.Y(n16),
	.B(P_data[2]),
	.A(n37), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U19 (
	.Y(n12),
	.A(P_data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U20 (
	.Y(n37),
	.A(P_data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U21 (
	.Y(n38),
	.A(P_data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U22 (
	.Y(n13),
	.A(P_data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U23 (
	.Y(n36),
	.A(P_data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U24 (
	.Y(n35),
	.A(P_data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U25 (
	.Y(n39),
	.A(P_data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U26 (
	.Y(N8),
	.B(prescale[5]),
	.A(\add_17/carry[4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U36 (
	.Y(N7),
	.B(\add_17/carry[4] ),
	.A(prescale[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U37 (
	.Y(\add_17/carry[4] ),
	.B(prescale[4]),
	.A(\add_17/carry[3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U38 (
	.Y(N6),
	.B(\add_17/carry[3] ),
	.A(prescale[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U39 (
	.Y(\add_17/carry[3] ),
	.B(prescale[3]),
	.A(prescale[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U40 (
	.Y(N5),
	.B(prescale[2]),
	.A(prescale[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U41 (
	.Y(n1),
	.B(N3),
	.AN(edge_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U42 (
	.Y(n6),
	.B1(n1),
	.B0(edge_count[1]),
	.A1N(N4),
	.A0(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U43 (
	.Y(n2),
	.B(edge_count[0]),
	.AN(N3), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U44 (
	.Y(n4),
	.B1(n2),
	.B0(N4),
	.A1N(edge_count[1]),
	.A0(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U45 (
	.Y(n3),
	.B(edge_count[5]),
	.A(N8), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X1M U46 (
	.Y(n10),
	.C(n3),
	.B(n4),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U47 (
	.Y(n9),
	.B(edge_count[4]),
	.A(N7), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U48 (
	.Y(n8),
	.B(edge_count[2]),
	.A(N5), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U49 (
	.Y(n7),
	.B(edge_count[3]),
	.A(N6), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U50 (
	.Y(N9),
	.D(n7),
	.C(n8),
	.B(n9),
	.A(n10), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module parity_chk_test_1 (
	clk, 
	rst, 
	parity_bit, 
	disable_err, 
	par_chk_en, 
	sampled_bit, 
	par_err, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input clk;
   input rst;
   input parity_bit;
   input disable_err;
   input par_chk_en;
   input sampled_bit;
   output par_err;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n2;
   wire n4;
   wire n5;
   wire n7;
   wire n8;
   wire n1;

   // Module instantiations
   OAI32X1M U6 (
	.Y(n5),
	.B1(n7),
	.B0(n4),
	.A2(disable_err),
	.A1(par_chk_en),
	.A0(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U7 (
	.Y(n4),
	.B(parity_bit),
	.A(sampled_bit), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U8 (
	.Y(n7),
	.A(par_chk_en), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M par_err_reg (
	.SI(parity_bit),
	.SE(test_se),
	.RN(rst),
	.QN(n2),
	.Q(n8),
	.D(n5),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U3 (
	.Y(n1),
	.A(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX12M U4 (
	.Y(par_err),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U5 (
	.Y(test_so),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module strt_chk (
	sampled_bit, 
	strt_chk_en, 
	strt_err, 
	VDD, 
	VSS);
   input sampled_bit;
   input strt_chk_en;
   output strt_err;
   inout VDD;
   inout VSS;

   // Module instantiations
   AND2X2M U2 (
	.Y(strt_err),
	.B(sampled_bit),
	.A(strt_chk_en), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module stp_chk (
	sampled_bit, 
	stp_chk_en, 
	stp_chk_err, 
	VDD, 
	VSS);
   input sampled_bit;
   input stp_chk_en;
   output stp_chk_err;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n2;

   // Module instantiations
   BUFX10M U2 (
	.Y(stp_chk_err),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U3 (
	.Y(n2),
	.B(sampled_bit),
	.AN(stp_chk_en), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module UART_TX_test_1 (
	clk, 
	rst, 
	data, 
	data_valid, 
	parity_enable, 
	parity_type, 
	TX_OUT, 
	busy, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN2_rst_from_sync2, 
	tx_clock__L3_N2, 
	tx_clock__L3_N3, 
	VDD, 
	VSS);
   input clk;
   input rst;
   input [7:0] data;
   input data_valid;
   input parity_enable;
   input parity_type;
   output TX_OUT;
   output busy;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN2_rst_from_sync2;
   input tx_clock__L3_N2;
   input tx_clock__L3_N3;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n11;
   wire serial_done;
   wire serial_enable;
   wire serial_data;
   wire parity_bit;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n13;
   wire [3:0] mux_select;

   // Module instantiations
   AOI21BX2M U3 (
	.Y(n11),
	.B0N(n5),
	.A1(n4),
	.A0(serial_data), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX12M U4 (
	.Y(TX_OUT),
	.A(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI32XLM U5 (
	.Y(n5),
	.B1(n7),
	.B0(parity_bit),
	.A2(n9),
	.A1(n6),
	.A0(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U6 (
	.Y(n10),
	.A(mux_select[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4BX1M U7 (
	.Y(n7),
	.D(mux_select[3]),
	.C(mux_select[1]),
	.B(mux_select[0]),
	.AN(mux_select[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U8 (
	.Y(n4),
	.D(mux_select[3]),
	.C(mux_select[2]),
	.B(mux_select[0]),
	.A(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BBX1M U9 (
	.Y(n6),
	.D(n10),
	.C(mux_select[0]),
	.BN(mux_select[3]),
	.AN(mux_select[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U12 (
	.Y(n8),
	.A(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U13 (
	.Y(n9),
	.A(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   FSM_test_1 controller (
	.clk(clk),
	.rst(rst),
	.data_valid(data_valid),
	.ser_done(serial_done),
	.parity_enable(parity_enable),
	.busy(busy),
	.ser_EN(serial_enable),
	.mux_sel({ mux_select[3],
		mux_select[2],
		mux_select[1],
		mux_select[0] }),
	.test_si(test_si),
	.test_so(n13),
	.test_se(test_se),
	.FE_OFN2_rst_from_sync2(FE_OFN2_rst_from_sync2),
	.tx_clock__L3_N3(tx_clock__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   serializer_test_1 ser (
	.clk(tx_clock__L3_N2),
	.rst(rst),
	.ser_EN(serial_enable),
	.dataValid(data_valid),
	.busy(busy),
	.data({ data[7],
		data[6],
		data[5],
		data[4],
		data[3],
		data[2],
		data[1],
		data[0] }),
	.ser_done(serial_done),
	.ser_data(serial_data),
	.test_si(parity_bit),
	.test_so(test_so),
	.test_se(test_se),
	.tx_clock__L3_N3(tx_clock__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   parityCalc_test_1 parity (
	.clk(clk),
	.rst(rst),
	.data({ data[7],
		data[6],
		data[5],
		data[4],
		data[3],
		data[2],
		data[1],
		data[0] }),
	.busy(busy),
	.data_valid(data_valid),
	.parity_type(parity_type),
	.parity_enable(parity_enable),
	.parity_bit(parity_bit),
	.test_si(n13),
	.test_se(test_se),
	.FE_OFN2_rst_from_sync2(FE_OFN2_rst_from_sync2),
	.tx_clock__L3_N2(tx_clock__L3_N2),
	.tx_clock__L3_N3(tx_clock__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module FSM_test_1 (
	clk, 
	rst, 
	data_valid, 
	ser_done, 
	parity_enable, 
	busy, 
	ser_EN, 
	mux_sel, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN2_rst_from_sync2, 
	tx_clock__L3_N3, 
	VDD, 
	VSS);
   input clk;
   input rst;
   input data_valid;
   input ser_done;
   input parity_enable;
   output busy;
   output ser_EN;
   output [3:0] mux_sel;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN2_rst_from_sync2;
   input tx_clock__L3_N3;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire [2:0] current_state;
   wire [2:0] next_state;

   assign test_so = current_state[2] ;

   // Module instantiations
   SDFFRQX2M \current_state_reg[2]  (
	.SI(current_state[1]),
	.SE(test_se),
	.RN(rst),
	.Q(current_state[2]),
	.D(next_state[2]),
	.CK(tx_clock__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[1]  (
	.SI(n14),
	.SE(test_se),
	.RN(FE_OFN2_rst_from_sync2),
	.Q(current_state[1]),
	.D(next_state[1]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U7 (
	.Y(busy),
	.B(n9),
	.A(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U8 (
	.Y(mux_sel[0]),
	.B(current_state[1]),
	.A(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U9 (
	.Y(mux_sel[2]),
	.B(current_state[2]),
	.A(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U10 (
	.Y(mux_sel[3]),
	.B(n8),
	.AN(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI31X1M U11 (
	.Y(next_state[2]),
	.B0(n12),
	.A2(current_state[2]),
	.A1(parity_enable),
	.A0(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U12 (
	.Y(n7),
	.B(current_state[1]),
	.A(ser_done), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U13 (
	.Y(n12),
	.A(mux_sel[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U14 (
	.Y(n8),
	.B(n6),
	.A(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X2M U15 (
	.Y(next_state[0]),
	.C0(n13),
	.B0(n10),
	.A1(n9),
	.A0(ser_done), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U16 (
	.Y(n13),
	.A(mux_sel[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U17 (
	.Y(n10),
	.B0(data_valid),
	.A1(mux_sel[3]),
	.A0(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U18 (
	.Y(n11),
	.B(current_state[1]),
	.A(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U19 (
	.Y(n9),
	.B(n6),
	.A(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U20 (
	.Y(next_state[1]),
	.B0(current_state[2]),
	.A1(n6),
	.A0(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U21 (
	.Y(mux_sel[1]),
	.A(ser_EN), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3BX2M U22 (
	.Y(ser_EN),
	.C(current_state[2]),
	.B(n6),
	.AN(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \current_state_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(FE_OFN2_rst_from_sync2),
	.QN(n6),
	.Q(n14),
	.D(next_state[0]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module serializer_test_1 (
	clk, 
	rst, 
	ser_EN, 
	dataValid, 
	busy, 
	data, 
	ser_done, 
	ser_data, 
	test_si, 
	test_so, 
	test_se, 
	tx_clock__L3_N3, 
	VDD, 
	VSS);
   input clk;
   input rst;
   input ser_EN;
   input dataValid;
   input busy;
   input [7:0] data;
   output ser_done;
   output ser_data;
   input test_si;
   output test_so;
   input test_se;
   input tx_clock__L3_N3;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N23;
   wire N24;
   wire N25;
   wire N27;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n12;
   wire n13;
   wire n14;
   wire [7:1] data_reg;
   wire [2:0] count;

   assign test_so = data_reg[7] ;
   assign ser_done = N27 ;

   // Module instantiations
   SDFFRQX2M \data_reg_reg[0]  (
	.SI(n13),
	.SE(test_se),
	.RN(rst),
	.Q(ser_data),
	.D(n27),
	.CK(tx_clock__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \data_reg_reg[6]  (
	.SI(data_reg[5]),
	.SE(test_se),
	.RN(rst),
	.Q(data_reg[6]),
	.D(n29),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \data_reg_reg[5]  (
	.SI(data_reg[4]),
	.SE(test_se),
	.RN(rst),
	.Q(data_reg[5]),
	.D(n30),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \data_reg_reg[4]  (
	.SI(data_reg[3]),
	.SE(test_se),
	.RN(rst),
	.Q(data_reg[4]),
	.D(n31),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \data_reg_reg[3]  (
	.SI(data_reg[2]),
	.SE(test_se),
	.RN(rst),
	.Q(data_reg[3]),
	.D(n32),
	.CK(tx_clock__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \data_reg_reg[2]  (
	.SI(data_reg[1]),
	.SE(test_se),
	.RN(rst),
	.Q(data_reg[2]),
	.D(n33),
	.CK(tx_clock__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \data_reg_reg[1]  (
	.SI(ser_data),
	.SE(test_se),
	.RN(rst),
	.Q(data_reg[1]),
	.D(n34),
	.CK(tx_clock__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \data_reg_reg[7]  (
	.SI(data_reg[6]),
	.SE(test_se),
	.RN(rst),
	.Q(data_reg[7]),
	.D(n28),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \count_reg[1]  (
	.SI(count[0]),
	.SE(test_se),
	.RN(rst),
	.Q(count[1]),
	.D(N24),
	.CK(tx_clock__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \count_reg[2]  (
	.SI(n12),
	.SE(test_se),
	.RN(rst),
	.Q(count[2]),
	.D(N25),
	.CK(tx_clock__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \count_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(rst),
	.Q(count[0]),
	.D(N23),
	.CK(tx_clock__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U14 (
	.Y(n18),
	.B(busy),
	.AN(dataValid), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U15 (
	.Y(n17),
	.B(n18),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U16 (
	.Y(n14),
	.A(ser_EN), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U17 (
	.Y(n15),
	.B(n17),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U18 (
	.Y(n27),
	.B0(n16),
	.A1N(n15),
	.A0N(ser_data), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U19 (
	.Y(n16),
	.B1(n18),
	.B0(data[0]),
	.A1(n17),
	.A0(data_reg[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U20 (
	.Y(n34),
	.B0(n24),
	.A1N(n15),
	.A0N(data_reg[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U21 (
	.Y(n24),
	.B1(n18),
	.B0(data[1]),
	.A1(n17),
	.A0(data_reg[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U22 (
	.Y(n33),
	.B0(n23),
	.A1N(data_reg[2]),
	.A0N(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U23 (
	.Y(n23),
	.B1(n18),
	.B0(data[2]),
	.A1(n17),
	.A0(data_reg[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U24 (
	.Y(n32),
	.B0(n22),
	.A1N(data_reg[3]),
	.A0N(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U25 (
	.Y(n22),
	.B1(n18),
	.B0(data[3]),
	.A1(n17),
	.A0(data_reg[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U26 (
	.Y(n31),
	.B0(n21),
	.A1N(data_reg[4]),
	.A0N(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U27 (
	.Y(n21),
	.B1(n18),
	.B0(data[4]),
	.A1(n17),
	.A0(data_reg[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U28 (
	.Y(n30),
	.B0(n20),
	.A1N(data_reg[5]),
	.A0N(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U29 (
	.Y(n20),
	.B1(n18),
	.B0(data[5]),
	.A1(n17),
	.A0(data_reg[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U30 (
	.Y(n29),
	.B0(n19),
	.A1N(data_reg[6]),
	.A0N(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U31 (
	.Y(n19),
	.B1(n18),
	.B0(data[6]),
	.A1(n17),
	.A0(data_reg[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U32 (
	.Y(n28),
	.B1(n18),
	.B0(data[7]),
	.A1(data_reg[7]),
	.A0(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X2M U33 (
	.Y(N27),
	.C(count[1]),
	.B(count[2]),
	.A(count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U34 (
	.Y(N25),
	.B1(n14),
	.B0(n25),
	.A1N(N23),
	.A0N(count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI32X1M U35 (
	.Y(n25),
	.B1(n12),
	.B0(count[2]),
	.A2(count[1]),
	.A1(n13),
	.A0(count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U36 (
	.Y(n13),
	.A(count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U37 (
	.Y(N23),
	.B(count[0]),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U38 (
	.Y(N24),
	.B(n14),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U39 (
	.Y(n26),
	.B(n12),
	.A(count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U40 (
	.Y(n12),
	.A(count[1]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module parityCalc_test_1 (
	clk, 
	rst, 
	data, 
	busy, 
	data_valid, 
	parity_type, 
	parity_enable, 
	parity_bit, 
	test_si, 
	test_se, 
	FE_OFN2_rst_from_sync2, 
	tx_clock__L3_N2, 
	tx_clock__L3_N3, 
	VDD, 
	VSS);
   input clk;
   input rst;
   input [7:0] data;
   input busy;
   input data_valid;
   input parity_type;
   input parity_enable;
   output parity_bit;
   input test_si;
   input test_se;
   input FE_OFN2_rst_from_sync2;
   input tx_clock__L3_N2;
   input tx_clock__L3_N3;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n1;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n9;
   wire n11;
   wire n13;
   wire n15;
   wire n17;
   wire n19;
   wire n21;
   wire n23;
   wire n25;
   wire n2;
   wire [7:0] DATA_reg;

   // Module instantiations
   SDFFRQX2M parity_bit_reg (
	.SI(DATA_reg[7]),
	.SE(test_se),
	.RN(rst),
	.Q(parity_bit),
	.D(n9),
	.CK(tx_clock__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \DATA_reg_reg[5]  (
	.SI(DATA_reg[4]),
	.SE(test_se),
	.RN(FE_OFN2_rst_from_sync2),
	.Q(DATA_reg[5]),
	.D(n21),
	.CK(tx_clock__L3_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \DATA_reg_reg[1]  (
	.SI(DATA_reg[0]),
	.SE(test_se),
	.RN(FE_OFN2_rst_from_sync2),
	.Q(DATA_reg[1]),
	.D(n13),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \DATA_reg_reg[4]  (
	.SI(DATA_reg[3]),
	.SE(test_se),
	.RN(FE_OFN2_rst_from_sync2),
	.Q(DATA_reg[4]),
	.D(n19),
	.CK(tx_clock__L3_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \DATA_reg_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(FE_OFN2_rst_from_sync2),
	.Q(DATA_reg[0]),
	.D(n11),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \DATA_reg_reg[2]  (
	.SI(DATA_reg[1]),
	.SE(test_se),
	.RN(FE_OFN2_rst_from_sync2),
	.Q(DATA_reg[2]),
	.D(n15),
	.CK(tx_clock__L3_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \DATA_reg_reg[3]  (
	.SI(DATA_reg[2]),
	.SE(test_se),
	.RN(FE_OFN2_rst_from_sync2),
	.Q(DATA_reg[3]),
	.D(n17),
	.CK(tx_clock__L3_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \DATA_reg_reg[6]  (
	.SI(DATA_reg[5]),
	.SE(test_se),
	.RN(rst),
	.Q(DATA_reg[6]),
	.D(n23),
	.CK(tx_clock__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \DATA_reg_reg[7]  (
	.SI(DATA_reg[6]),
	.SE(test_se),
	.RN(rst),
	.Q(DATA_reg[7]),
	.D(n25),
	.CK(tx_clock__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U2 (
	.Y(n7),
	.B(busy),
	.AN(data_valid), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U3 (
	.Y(n5),
	.B(DATA_reg[3]),
	.A(DATA_reg[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U4 (
	.Y(n3),
	.C(n6),
	.B(DATA_reg[4]),
	.A(DATA_reg[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U5 (
	.Y(n6),
	.B(DATA_reg[6]),
	.A(DATA_reg[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U6 (
	.Y(n9),
	.B1(n2),
	.B0(n1),
	.A1N(n2),
	.A0N(parity_bit), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U7 (
	.Y(n2),
	.A(parity_enable), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U8 (
	.Y(n1),
	.C(n4),
	.B(parity_type),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U9 (
	.Y(n4),
	.C(n5),
	.B(DATA_reg[0]),
	.A(DATA_reg[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U10 (
	.Y(n11),
	.B1(n7),
	.B0(data[0]),
	.A1N(n7),
	.A0(DATA_reg[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U11 (
	.Y(n13),
	.B1(n7),
	.B0(data[1]),
	.A1N(n7),
	.A0(DATA_reg[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U12 (
	.Y(n15),
	.B1(n7),
	.B0(data[2]),
	.A1N(n7),
	.A0(DATA_reg[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U13 (
	.Y(n17),
	.B1(n7),
	.B0(data[3]),
	.A1N(n7),
	.A0(DATA_reg[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U14 (
	.Y(n19),
	.B1(n7),
	.B0(data[4]),
	.A1N(n7),
	.A0(DATA_reg[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U15 (
	.Y(n21),
	.B1(n7),
	.B0(data[5]),
	.A1N(n7),
	.A0(DATA_reg[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U16 (
	.Y(n23),
	.B1(n7),
	.B0(data[6]),
	.A1N(n7),
	.A0(DATA_reg[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U17 (
	.Y(n25),
	.B1(n7),
	.B0(data[7]),
	.A1N(n7),
	.A0(DATA_reg[7]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module DATA_SYNC_test_1 (
	unsync_bus, 
	bus_enable, 
	CLK, 
	RST, 
	sync_bus, 
	enable_pulse, 
	test_si2, 
	test_si1, 
	test_se, 
	ref_clock__L5_N1, 
	VDD, 
	VSS);
   input [7:0] unsync_bus;
   input bus_enable;
   input CLK;
   input RST;
   output [7:0] sync_bus;
   output enable_pulse;
   input test_si2;
   input test_si1;
   input test_se;
   input ref_clock__L5_N1;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN9_SI_1_;
   wire FE_PHN8_SI_1_;
   wire ex_enable;
   wire enable;
   wire exx_en;
   wire n1;
   wire n3;
   wire n5;
   wire n7;
   wire n9;
   wire n11;
   wire n13;
   wire n15;
   wire n17;
   wire n22;

   // Module instantiations
   DLY4X1M FE_PHC9_SI_1_ (
	.Y(FE_PHN9_SI_1_),
	.A(FE_PHN8_SI_1_), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC8_SI_1_ (
	.Y(FE_PHN8_SI_1_),
	.A(test_si2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M exx_en_reg (
	.SI(ex_enable),
	.SE(test_se),
	.RN(RST),
	.Q(exx_en),
	.D(ex_enable),
	.CK(ref_clock__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M ex_enable_reg (
	.SI(enable),
	.SE(test_se),
	.RN(RST),
	.Q(ex_enable),
	.D(enable),
	.CK(ref_clock__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M enable_pulse_reg (
	.SI(test_si1),
	.SE(test_se),
	.RN(RST),
	.Q(enable_pulse),
	.D(n22),
	.CK(ref_clock__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[7]  (
	.SI(sync_bus[6]),
	.SE(test_se),
	.RN(RST),
	.Q(sync_bus[7]),
	.D(n3),
	.CK(ref_clock__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[3]  (
	.SI(sync_bus[2]),
	.SE(test_se),
	.RN(RST),
	.Q(sync_bus[3]),
	.D(n11),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[6]  (
	.SI(sync_bus[5]),
	.SE(test_se),
	.RN(RST),
	.Q(sync_bus[6]),
	.D(n5),
	.CK(ref_clock__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[5]  (
	.SI(sync_bus[4]),
	.SE(test_se),
	.RN(RST),
	.Q(sync_bus[5]),
	.D(n7),
	.CK(ref_clock__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX4M \sync_bus_reg[1]  (
	.SI(sync_bus[0]),
	.SE(test_se),
	.RN(RST),
	.Q(sync_bus[1]),
	.D(n15),
	.CK(ref_clock__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[2]  (
	.SI(FE_PHN9_SI_1_),
	.SE(test_se),
	.RN(RST),
	.Q(sync_bus[2]),
	.D(n13),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[4]  (
	.SI(sync_bus[3]),
	.SE(test_se),
	.RN(RST),
	.Q(sync_bus[4]),
	.D(n9),
	.CK(ref_clock__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[0]  (
	.SI(exx_en),
	.SE(test_se),
	.RN(RST),
	.Q(sync_bus[0]),
	.D(n17),
	.CK(ref_clock__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M enable_reg (
	.SI(enable_pulse),
	.SE(test_se),
	.RN(RST),
	.Q(enable),
	.D(bus_enable),
	.CK(ref_clock__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U3 (
	.Y(n22),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U4 (
	.Y(n1),
	.B(ex_enable),
	.AN(exx_en), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U5 (
	.Y(n3),
	.B1(n1),
	.B0(sync_bus[7]),
	.A1(n22),
	.A0(unsync_bus[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U6 (
	.Y(n5),
	.B1(n1),
	.B0(sync_bus[6]),
	.A1(n22),
	.A0(unsync_bus[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U7 (
	.Y(n7),
	.B1(n1),
	.B0(sync_bus[5]),
	.A1(n22),
	.A0(unsync_bus[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U8 (
	.Y(n9),
	.B1(n1),
	.B0(sync_bus[4]),
	.A1(n22),
	.A0(unsync_bus[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U9 (
	.Y(n11),
	.B1(n1),
	.B0(sync_bus[3]),
	.A1(n22),
	.A0(unsync_bus[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U10 (
	.Y(n13),
	.B1(n1),
	.B0(sync_bus[2]),
	.A1(n22),
	.A0(unsync_bus[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U11 (
	.Y(n15),
	.B1(n1),
	.B0(sync_bus[1]),
	.A1(n22),
	.A0(unsync_bus[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U12 (
	.Y(n17),
	.B1(n1),
	.B0(sync_bus[0]),
	.A1(n22),
	.A0(unsync_bus[0]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module CLK_GATE (
	CLK_EN, 
	CLK, 
	test_en, 
	GATED_CLK, 
	VDD, 
	VSS);
   input CLK_EN;
   input CLK;
   input test_en;
   output GATED_CLK;
   inout VDD;
   inout VSS;

   // Internal wires
   wire _0_net_;

   // Module instantiations
   TLATNCAX16M u0 (
	.ECK(GATED_CLK),
	.E(_0_net_),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U1 (
	.Y(_0_net_),
	.B(test_en),
	.A(CLK_EN), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module PULSE_GEN_test_0 (
	CLK, 
	RST, 
	LVL_SIG, 
	PULSE_SIG, 
	test_si, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input LVL_SIG;
   output PULSE_SIG;
   input test_si;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire internal;
   wire pulse;

   assign test_so = internal ;

   // Module instantiations
   SDFFRQX2M internal_reg (
	.SI(PULSE_SIG),
	.SE(test_se),
	.RN(RST),
	.Q(internal),
	.D(LVL_SIG),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M PULSE_SIG_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(PULSE_SIG),
	.D(pulse),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U5 (
	.Y(pulse),
	.B(internal),
	.AN(LVL_SIG), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module PULSE_GEN_test_1 (
	CLK, 
	RST, 
	LVL_SIG, 
	PULSE_SIG, 
	test_si, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input LVL_SIG;
   output PULSE_SIG;
   input test_si;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire internal;
   wire pulse;

   assign test_so = internal ;

   // Module instantiations
   SDFFRQX2M internal_reg (
	.SI(PULSE_SIG),
	.SE(test_se),
	.RN(RST),
	.Q(internal),
	.D(LVL_SIG),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M PULSE_SIG_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(PULSE_SIG),
	.D(pulse),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U5 (
	.Y(pulse),
	.B(internal),
	.AN(LVL_SIG), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module PULSE_SAMEZERO_GEN_test_1 (
	CLK, 
	RST, 
	busyFall, 
	empty, 
	PULSE_SIG, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input busyFall;
   input empty;
   output PULSE_SIG;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N4;

   // Module instantiations
   SDFFRQX4M PULSE_SIG_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(PULSE_SIG),
	.D(N4),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U4 (
	.Y(N4),
	.B(busyFall),
	.AN(empty), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module PULSE_NEG_GEN_test_1 (
	CLK, 
	RST, 
	LVL_SIG, 
	PULSE_SIG, 
	test_si, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input LVL_SIG;
   output PULSE_SIG;
   input test_si;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire internal;
   wire n3;

   assign test_so = internal ;

   // Module instantiations
   SDFFRQX2M internal_reg (
	.SI(PULSE_SIG),
	.SE(test_se),
	.RN(RST),
	.Q(internal),
	.D(LVL_SIG),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M PULSE_SIG_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(PULSE_SIG),
	.D(n3),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U5 (
	.Y(n3),
	.B(LVL_SIG),
	.AN(internal), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ClkDiv_test_0 (
	i_ref_clk, 
	i_rst_n, 
	i_clk_en, 
	i_div_ratio, 
	o_div_clk, 
	test_si, 
	test_so, 
	test_se, 
	n12__Exclude_0_NET, 
	uart_clock__L3_N0, 
	uart_clock__L7_N0, 
	VDD, 
	VSS);
   input i_ref_clk;
   input i_rst_n;
   input i_clk_en;
   input [7:0] i_div_ratio;
   output o_div_clk;
   input test_si;
   output test_so;
   input test_se;
   input n12__Exclude_0_NET;
   input uart_clock__L3_N0;
   input uart_clock__L7_N0;
   inout VDD;
   inout VSS;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire N1;
   wire o_div_clk_;
   wire flag;
   wire N7;
   wire N11;
   wire N12;
   wire N13;
   wire N14;
   wire N15;
   wire N16;
   wire N17;
   wire N18;
   wire N19;
   wire N26;
   wire N27;
   wire N28;
   wire N29;
   wire N30;
   wire N31;
   wire N32;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n1;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n17;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire [6:0] count;

//   assign test_so = o_div_clk_ ;

   // Module instantiations
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSQX2M flag_reg (
	.SN(i_rst_n),
	.SI(count[6]),
	.SE(test_se),
	.Q(flag),
	.D(n36),
	.CK(i_ref_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M o_div_clk__reg (
	.SI(flag),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(test_so),
	.D(n28),
	.CK(uart_clock__L3_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \count_reg[6]  (
	.SI(count[5]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(count[6]),
	.D(n35),
	.CK(i_ref_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSQX2M \count_reg[0]  (
	.SN(i_rst_n),
	.SI(test_si),
	.SE(test_se),
	.Q(count[0]),
	.D(n34),
	.CK(i_ref_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \count_reg[3]  (
	.SI(count[2]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(count[3]),
	.D(n31),
	.CK(i_ref_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \count_reg[2]  (
	.SI(count[1]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(count[2]),
	.D(n32),
	.CK(i_ref_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \count_reg[5]  (
	.SI(count[4]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(count[5]),
	.D(n29),
	.CK(i_ref_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \count_reg[4]  (
	.SI(count[3]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(count[4]),
	.D(n30),
	.CK(i_ref_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \count_reg[1]  (
	.SI(count[0]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(count[1]),
	.D(n33),
	.CK(i_ref_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U5 (
	.Y(n19),
	.B(n20),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U7 (
	.Y(n25),
	.C(N7),
	.B(n51),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   AND4X2M U11 (
	.Y(n20),
	.D(n25),
	.C(n24),
	.B(n23),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U16 (
	.Y(n18),
	.C(n23),
	.B(n25),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U17 (
	.Y(N1),
	.B(n26),
	.A(n51), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U18 (
	.Y(n24),
	.D(n22),
	.C(N7),
	.B(flag),
	.A(i_div_ratio[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BX1M U19 (
	.Y(n23),
	.D(n22),
	.C(i_div_ratio[0]),
	.B(N19),
	.AN(flag), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U20 (
	.Y(n34),
	.B(n21),
	.AN(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U21 (
	.Y(n21),
	.B1(n19),
	.B0(count[0]),
	.A1(n20),
	.A0(N26), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U22 (
	.Y(n33),
	.B1(n20),
	.B0(N27),
	.A1(n19),
	.A0(count[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U23 (
	.Y(n32),
	.B1(n20),
	.B0(N28),
	.A1(n19),
	.A0(count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U24 (
	.Y(n31),
	.B1(n20),
	.B0(N29),
	.A1(n19),
	.A0(count[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U25 (
	.Y(n30),
	.B1(n20),
	.B0(N30),
	.A1(n19),
	.A0(count[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U26 (
	.Y(n29),
	.B1(n20),
	.B0(N31),
	.A1(n19),
	.A0(count[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U27 (
	.Y(n35),
	.B1(n20),
	.B0(N32),
	.A1(n19),
	.A0(count[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U28 (
	.Y(n36),
	.B0(n23),
	.A1N(flag),
	.A0N(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U29 (
	.Y(n22),
	.B(n26),
	.A(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   OR4X1M U30 (
	.Y(n26),
	.D(n27),
	.C(i_div_ratio[1]),
	.B(i_div_ratio[2]),
	.A(i_div_ratio[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR4X1M U31 (
	.Y(n27),
	.D(i_div_ratio[6]),
	.C(i_div_ratio[7]),
	.B(i_div_ratio[4]),
	.A(i_div_ratio[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U32 (
	.Y(n28),
	.B(n12__Exclude_0_NET),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U33 (
	.Y(n51),
	.A(i_div_ratio[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U34 (
	.Y(o_div_clk),
	.S0(N1),
	.B(uart_clock__L7_N0),
	.A(test_so), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U35 (
	.Y(n7),
	.B(count[3]),
	.A(i_div_ratio[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U36 (
	.Y(n6),
	.B(count[2]),
	.A(i_div_ratio[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U37 (
	.Y(n1),
	.B(count[0]),
	.AN(i_div_ratio[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U38 (
	.Y(n5),
	.B1(n1),
	.B0(i_div_ratio[2]),
	.A1N(count[1]),
	.A0(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U39 (
	.Y(n3),
	.B(i_div_ratio[1]),
	.AN(count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U40 (
	.Y(n4),
	.B1(n3),
	.B0(count[1]),
	.A1N(i_div_ratio[2]),
	.A0(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X1M U41 (
	.Y(n39),
	.D(n4),
	.C(n5),
	.B(n6),
	.A(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U42 (
	.Y(n38),
	.B(count[6]),
	.A(i_div_ratio[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U43 (
	.Y(n37),
	.B(count[4]),
	.A(i_div_ratio[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U44 (
	.Y(n17),
	.B(count[5]),
	.A(i_div_ratio[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U45 (
	.Y(N7),
	.D(n17),
	.C(n37),
	.B(n38),
	.A(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U46 (
	.Y(n40),
	.B(count[0]),
	.AN(N11), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U47 (
	.Y(n44),
	.B1(n40),
	.B0(N12),
	.A1N(count[1]),
	.A0(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U48 (
	.Y(n43),
	.B(count[2]),
	.A(N13), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U49 (
	.Y(n41),
	.B(N11),
	.AN(count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U50 (
	.Y(n42),
	.B1(n41),
	.B0(count[1]),
	.A1N(N12),
	.A0(n41), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BX1M U51 (
	.Y(n50),
	.D(n42),
	.C(n43),
	.B(n44),
	.AN(N18), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U52 (
	.Y(n48),
	.B(count[6]),
	.A(N17), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U53 (
	.Y(n47),
	.B(count[5]),
	.A(N16), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U54 (
	.Y(n46),
	.B(count[4]),
	.A(N15), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U55 (
	.Y(n45),
	.B(count[3]),
	.A(N14), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X1M U56 (
	.Y(n49),
	.D(n45),
	.C(n46),
	.B(n47),
	.A(n48), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U57 (
	.Y(N19),
	.B(n49),
	.A(n50), 
	.VDD(VDD), 
	.VSS(VSS));
   ClkDiv_0_DW01_inc_0 add_36 (
	.A({ count[6],
		count[5],
		count[4],
		count[3],
		count[2],
		count[1],
		count[0] }),
	.SUM({ N32,
		N31,
		N30,
		N29,
		N28,
		N27,
		N26 }), 
	.VDD(VDD), 
	.VSS(VSS));
   ClkDiv_0_DW01_inc_1 add_30 (
	.A({ 1'b0,
		i_div_ratio[7],
		i_div_ratio[6],
		i_div_ratio[5],
		i_div_ratio[4],
		i_div_ratio[3],
		i_div_ratio[2],
		i_div_ratio[1] }),
	.SUM({ N18,
		N17,
		N16,
		N15,
		N14,
		N13,
		N12,
		N11 }), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ClkDiv_0_DW01_inc_0 (
	A, 
	SUM, 
	VDD, 
	VSS);
   input [6:0] A;
   output [6:0] SUM;
   inout VDD;
   inout VSS;

   // Internal wires
   wire [6:2] carry;

   // Module instantiations
   ADDHX1M U1_1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.B(carry[5]),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.B(carry[4]),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.B(carry[3]),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.B(carry[2]),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.B(A[0]),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U1 (
	.Y(SUM[6]),
	.B(A[6]),
	.A(carry[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U2 (
	.Y(SUM[0]),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ClkDiv_0_DW01_inc_1 (
	A, 
	SUM, 
	VDD, 
	VSS);
   input [7:0] A;
   output [7:0] SUM;
   inout VDD;
   inout VSS;

   // Internal wires
   wire [7:2] carry;

   // Module instantiations
   ADDHX1M U1_1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.B(carry[4]),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.B(carry[3]),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.B(carry[2]),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.B(A[0]),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.B(carry[5]),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_6 (
	.S(SUM[6]),
	.CO(SUM[7]),
	.B(carry[6]),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U1 (
	.Y(SUM[0]),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ClkDiv_test_1 (
	i_ref_clk, 
	i_rst_n, 
	i_clk_en, 
	i_div_ratio, 
	o_div_clk, 
	test_si, 
	test_so, 
	test_se, 
	n11__Exclude_0_NET, 
	uart_clock__L3_N1, 
	uart_clock__L7_N1, 
	VDD, 
	VSS);
   input i_ref_clk;
   input i_rst_n;
   input i_clk_en;
   input [7:0] i_div_ratio;
   output o_div_clk;
   input test_si;
   output test_so;
   input test_se;
   input n11__Exclude_0_NET;
   input uart_clock__L3_N1;
   input uart_clock__L7_N1;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN17_n12__Exclude_0_NET;
   wire HTIE_LTIEHI_NET;
   wire LTIE_LTIELO_NET;
   wire N1;
   wire o_div_clk_;
   wire flag;
   wire N7;
   wire N11;
   wire N12;
   wire N13;
   wire N14;
   wire N15;
   wire N16;
   wire N17;
   wire N18;
   wire N19;
   wire N26;
   wire N27;
   wire N28;
   wire N29;
   wire N30;
   wire N31;
   wire N32;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n17;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire [6:0] count;

//   assign test_so = o_div_clk_ ;

   // Module instantiations
   DLY4X1M FE_PHC17_n12__Exclude_0_NET (
	.Y(FE_PHN17_n12__Exclude_0_NET),
	.A(test_si), 
	.VDD(VDD), 
	.VSS(VSS));
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   TIELOM LTIE_LTIELO (
	.Y(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M o_div_clk__reg (
	.SI(flag),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(test_so),
	.D(n61),
	.CK(uart_clock__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \count_reg[6]  (
	.SI(count[5]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(count[6]),
	.D(n54),
	.CK(i_ref_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSQX2M \count_reg[0]  (
	.SN(i_rst_n),
	.SI(FE_PHN17_n12__Exclude_0_NET),
	.SE(test_se),
	.Q(count[0]),
	.D(n55),
	.CK(i_ref_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \count_reg[3]  (
	.SI(count[2]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(count[3]),
	.D(n58),
	.CK(i_ref_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \count_reg[2]  (
	.SI(count[1]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(count[2]),
	.D(n57),
	.CK(i_ref_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \count_reg[5]  (
	.SI(count[4]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(count[5]),
	.D(n60),
	.CK(i_ref_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \count_reg[4]  (
	.SI(count[3]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(count[4]),
	.D(n59),
	.CK(i_ref_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \count_reg[1]  (
	.SI(count[0]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(count[1]),
	.D(n56),
	.CK(i_ref_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSQX1M flag_reg (
	.SN(i_rst_n),
	.SI(count[6]),
	.SE(test_se),
	.Q(flag),
	.D(n53),
	.CK(i_ref_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U7 (
	.Y(n70),
	.B(n69),
	.A(n71), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U11 (
	.Y(n64),
	.C(N7),
	.B(n52),
	.A(n67), 
	.VDD(VDD), 
	.VSS(VSS));
   AND4X2M U16 (
	.Y(n69),
	.D(n64),
	.C(n65),
	.B(n66),
	.A(n67), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U17 (
	.Y(n71),
	.C(n66),
	.B(n64),
	.A(n65), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U18 (
	.Y(n52),
	.A(i_div_ratio[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U19 (
	.Y(N1),
	.B(n63),
	.A(n52), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U20 (
	.Y(n65),
	.D(n67),
	.C(N7),
	.B(flag),
	.A(i_div_ratio[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U21 (
	.Y(n55),
	.B(n68),
	.AN(n71), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U22 (
	.Y(n68),
	.B1(n70),
	.B0(count[0]),
	.A1(n69),
	.A0(N26), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U23 (
	.Y(n56),
	.B1(n69),
	.B0(N27),
	.A1(n70),
	.A0(count[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U24 (
	.Y(n57),
	.B1(n69),
	.B0(N28),
	.A1(n70),
	.A0(count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U25 (
	.Y(n58),
	.B1(n69),
	.B0(N29),
	.A1(n70),
	.A0(count[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U26 (
	.Y(n59),
	.B1(n69),
	.B0(N30),
	.A1(n70),
	.A0(count[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U27 (
	.Y(n60),
	.B1(n69),
	.B0(N31),
	.A1(n70),
	.A0(count[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U28 (
	.Y(n54),
	.B1(n69),
	.B0(N32),
	.A1(n70),
	.A0(count[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BX1M U29 (
	.Y(n66),
	.D(n67),
	.C(i_div_ratio[0]),
	.B(N19),
	.AN(flag), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U30 (
	.Y(n53),
	.B0(n66),
	.A1N(flag),
	.A0N(n65), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U31 (
	.Y(n67),
	.B(n63),
	.A(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   OR4X1M U32 (
	.Y(n63),
	.D(n62),
	.C(i_div_ratio[1]),
	.B(i_div_ratio[2]),
	.A(i_div_ratio[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR4X1M U33 (
	.Y(n62),
	.D(LTIE_LTIELO_NET),
	.C(LTIE_LTIELO_NET),
	.B(LTIE_LTIELO_NET),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U34 (
	.Y(n61),
	.B(n11__Exclude_0_NET),
	.A(n71), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U35 (
	.Y(o_div_clk),
	.S0(N1),
	.B(uart_clock__L7_N1),
	.A(test_so), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U36 (
	.Y(n17),
	.B(count[3]),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U37 (
	.Y(n7),
	.B(count[2]),
	.A(i_div_ratio[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U38 (
	.Y(n3),
	.B(count[0]),
	.AN(i_div_ratio[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U39 (
	.Y(n6),
	.B1(n3),
	.B0(i_div_ratio[2]),
	.A1N(count[1]),
	.A0(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U40 (
	.Y(n4),
	.B(i_div_ratio[1]),
	.AN(count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U41 (
	.Y(n5),
	.B1(n4),
	.B0(count[1]),
	.A1N(i_div_ratio[2]),
	.A0(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X1M U42 (
	.Y(n40),
	.D(n5),
	.C(n6),
	.B(n7),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U43 (
	.Y(n39),
	.B(count[6]),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U44 (
	.Y(n38),
	.B(count[4]),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U45 (
	.Y(n37),
	.B(count[5]),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U46 (
	.Y(N7),
	.D(n37),
	.C(n38),
	.B(n39),
	.A(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U47 (
	.Y(n41),
	.B(count[0]),
	.AN(N11), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U48 (
	.Y(n45),
	.B1(n41),
	.B0(N12),
	.A1N(count[1]),
	.A0(n41), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U49 (
	.Y(n44),
	.B(count[2]),
	.A(N13), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U50 (
	.Y(n42),
	.B(N11),
	.AN(count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U51 (
	.Y(n43),
	.B1(n42),
	.B0(count[1]),
	.A1N(N12),
	.A0(n42), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BX1M U52 (
	.Y(n51),
	.D(n43),
	.C(n44),
	.B(n45),
	.AN(N18), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U53 (
	.Y(n49),
	.B(count[6]),
	.A(N17), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U54 (
	.Y(n48),
	.B(count[5]),
	.A(N16), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U55 (
	.Y(n47),
	.B(count[4]),
	.A(N15), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U56 (
	.Y(n46),
	.B(count[3]),
	.A(N14), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X1M U57 (
	.Y(n50),
	.D(n46),
	.C(n47),
	.B(n48),
	.A(n49), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U58 (
	.Y(N19),
	.B(n50),
	.A(n51), 
	.VDD(VDD), 
	.VSS(VSS));
   ClkDiv_1_DW01_inc_0 add_36 (
	.A({ count[6],
		count[5],
		count[4],
		count[3],
		count[2],
		count[1],
		count[0] }),
	.SUM({ N32,
		N31,
		N30,
		N29,
		N28,
		N27,
		N26 }), 
	.VDD(VDD), 
	.VSS(VSS));
   ClkDiv_1_DW01_inc_1 add_30 (
	.A({ 1'b0,
		i_div_ratio[7],
		i_div_ratio[6],
		i_div_ratio[5],
		i_div_ratio[4],
		i_div_ratio[3],
		i_div_ratio[2],
		i_div_ratio[1] }),
	.SUM({ N18,
		N17,
		N16,
		N15,
		N14,
		N13,
		N12,
		N11 }), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ClkDiv_1_DW01_inc_0 (
	A, 
	SUM, 
	VDD, 
	VSS);
   input [6:0] A;
   output [6:0] SUM;
   inout VDD;
   inout VSS;

   // Internal wires
   wire [6:2] carry;

   // Module instantiations
   ADDHX1M U1_1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.B(carry[5]),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.B(carry[4]),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.B(carry[3]),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.B(carry[2]),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.B(A[0]),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U1 (
	.Y(SUM[6]),
	.B(A[6]),
	.A(carry[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U2 (
	.Y(SUM[0]),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ClkDiv_1_DW01_inc_1 (
	A, 
	SUM, 
	VDD, 
	VSS);
   input [7:0] A;
   output [7:0] SUM;
   inout VDD;
   inout VSS;

   // Internal wires
   wire LTIE_LTIELO_NET;
   wire [7:2] carry;

   // Module instantiations
   TIELOM LTIE_LTIELO (
	.Y(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_6 (
	.S(SUM[6]),
	.CO(SUM[7]),
	.B(carry[6]),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.B(carry[5]),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.B(carry[4]),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.B(carry[3]),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.B(carry[2]),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.B(A[0]),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U1 (
	.Y(SUM[0]),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module RST_SYNC_test_0 (
	CLK, 
	RST, 
	SYNC_RST, 
	test_si, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   output SYNC_RST;
   input test_si;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN16_n11__Exclude_0_NET;
   wire HTIE_LTIEHI_NET;
   wire internal;

   assign test_so = internal ;

   // Module instantiations
   DLY4X1M FE_PHC16_n11__Exclude_0_NET (
	.Y(FE_PHN16_n11__Exclude_0_NET),
	.A(test_si), 
	.VDD(VDD), 
	.VSS(VSS));
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M internal_reg (
	.SI(SYNC_RST),
	.SE(test_se),
	.RN(RST),
	.Q(internal),
	.D(HTIE_LTIEHI_NET),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX1M SYNC_RST_reg (
	.SI(FE_PHN16_n11__Exclude_0_NET),
	.SE(test_se),
	.RN(RST),
	.Q(SYNC_RST),
	.D(internal),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module RST_SYNC_test_1 (
	CLK, 
	RST, 
	SYNC_RST, 
	test_si, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   output SYNC_RST;
   input test_si;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire internal;

   assign test_so = internal ;

   // Module instantiations
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M internal_reg (
	.SI(SYNC_RST),
	.SE(test_se),
	.RN(RST),
	.Q(internal),
	.D(HTIE_LTIEHI_NET),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX1M SYNC_RST_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(SYNC_RST),
	.D(internal),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module custom_mux (
	selector, 
	div_ratio, 
	VDD, 
	VSS);
   input [5:0] selector;
   output [7:0] div_ratio;
   inout VDD;
   inout VSS;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n14;
   wire n15;
   wire n16;
   wire n17;

   // Module instantiations
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U11 (
	.Y(div_ratio[3]),
	.D(selector[4]),
	.C(selector[5]),
	.B(selector[3]),
	.A(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U12 (
	.Y(div_ratio[2]),
	.C(selector[0]),
	.B(selector[1]),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BX1M U13 (
	.Y(n6),
	.D(n14),
	.C(n15),
	.B(selector[3]),
	.AN(selector[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BX1M U14 (
	.Y(n7),
	.D(n14),
	.C(n15),
	.B(selector[4]),
	.AN(selector[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U15 (
	.Y(div_ratio[1]),
	.C(selector[0]),
	.B(selector[1]),
	.A(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U16 (
	.Y(n15),
	.A(selector[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U17 (
	.Y(n14),
	.A(selector[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U18 (
	.Y(n5),
	.C(selector[2]),
	.B(n16),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U19 (
	.Y(n16),
	.A(selector[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U20 (
	.Y(n17),
	.A(selector[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X2M U21 (
	.Y(div_ratio[0]),
	.C0(n16),
	.B0(n17),
	.A1(n9),
	.A0(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U22 (
	.Y(n8),
	.D(n15),
	.C(selector[3]),
	.B(selector[4]),
	.A(selector[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U23 (
	.Y(n9),
	.B(n6),
	.A(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U3 (
	.Y(div_ratio[4]),
	.A(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U5 (
	.Y(div_ratio[5]),
	.A(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U7 (
	.Y(div_ratio[6]),
	.A(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U9 (
	.Y(div_ratio[7]),
	.A(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SYS_TOP (
	REF_CLK, 
	UART_CLK, 
	RST, 
	RX_IN, 
	SI, 
	SE, 
	test_mode, 
	scan_clk, 
	scan_rst, 
	SO, 
	TX_OUT, 
	parity_error, 
	frame_error, 
	VDD, 
	VSS);
   input REF_CLK;
   input UART_CLK;
   input RST;
   input RX_IN;
   input [3:0] SI;
   input SE;
   input test_mode;
   input scan_clk;
   input scan_rst;
   output [3:0] SO;
   output TX_OUT;
   output parity_error;
   output frame_error;
   inout VDD;
   inout VSS;

   // Internal wires
   wire REF_CLK__L2_N0;
   wire REF_CLK__L1_N0;
   wire UART_CLK__L2_N0;
   wire UART_CLK__L1_N0;
   wire scan_clk__L12_N0;
   wire scan_clk__L11_N0;
   wire scan_clk__L10_N0;
   wire scan_clk__L9_N1;
   wire scan_clk__L9_N0;
   wire scan_clk__L8_N1;
   wire scan_clk__L8_N0;
   wire scan_clk__L7_N1;
   wire scan_clk__L7_N0;
   wire scan_clk__L6_N1;
   wire scan_clk__L6_N0;
   wire scan_clk__L5_N1;
   wire scan_clk__L5_N0;
   wire scan_clk__L4_N0;
   wire scan_clk__L3_N0;
   wire scan_clk__L2_N0;
   wire scan_clk__L1_N0;
   wire ref_clock__L5_N7;
   wire ref_clock__L5_N6;
   wire ref_clock__L5_N5;
   wire ref_clock__L5_N4;
   wire ref_clock__L5_N3;
   wire ref_clock__L5_N2;
   wire ref_clock__L5_N1;
   wire ref_clock__L5_N0;
   wire ref_clock__L4_N3;
   wire ref_clock__L4_N2;
   wire ref_clock__L4_N1;
   wire ref_clock__L4_N0;
   wire ref_clock__L3_N1;
   wire ref_clock__L3_N0;
   wire ref_clock__L2_N0;
   wire ref_clock__L1_N0;
   wire gated_clk__L3_N1;
   wire gated_clk__L3_N0;
   wire gated_clk__L2_N0;
   wire gated_clk__L1_N0;
   wire uart_clock__L12_N1;
   wire uart_clock__L12_N0;
   wire uart_clock__L11_N0;
   wire uart_clock__L10_N0;
   wire uart_clock__L9_N0;
   wire uart_clock__L8_N0;
   wire uart_clock__L7_N2;
   wire uart_clock__L7_N1;
   wire uart_clock__L7_N0;
   wire uart_clock__L6_N1;
   wire uart_clock__L6_N0;
   wire uart_clock__L5_N1;
   wire uart_clock__L5_N0;
   wire uart_clock__L4_N0;
   wire uart_clock__L3_N2;
   wire uart_clock__L3_N1;
   wire uart_clock__L3_N0;
   wire uart_clock__L2_N0;
   wire uart_clock__L1_N0;
   wire n12__Exclude_0_NET;
   wire n11__Exclude_0_NET;
   wire tx_clock__L3_N3;
   wire tx_clock__L3_N2;
   wire tx_clock__L3_N1;
   wire tx_clock__L3_N0;
   wire tx_clock__L2_N0;
   wire tx_clock__L1_N0;
   wire rx_clock__L3_N3;
   wire rx_clock__L3_N2;
   wire rx_clock__L3_N1;
   wire rx_clock__L3_N0;
   wire rx_clock__L2_N0;
   wire rx_clock__L1_N0;
   wire FE_OFN5_SE;
   wire FE_OFN2_rst_from_sync2;
   wire FE_OFN1_rst_from_sync1;
   wire FE_OFN0_rst_from_sync1;
   wire ref_clock;
   wire uart_clock;
   wire TX_CLK;
   wire tx_clock;
   wire RX_CLK;
   wire rx_clock;
   wire rst_to_sync;
   wire sync_rst1;
   wire rst_from_sync1;
   wire sync_rst2;
   wire rst_from_sync2;
   wire write_enable_reg;
   wire read_enable_reg;
   wire read_valid_reg;
   wire alu_enable;
   wire gated_clk;
   wire out_valid;
   wire rx_d_valid;
   wire full;
   wire tx_idle;
   wire clock_gate_enable;
   wire write_inc;
   wire read_inc;
   wire empty;
   wire rx_out_valid;
   wire vld;
   wire busy;
   wire pulsing_empty;
   wire n1;
   wire n2;
   wire n3;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n21;
   wire n22;
   wire n25;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire [7:0] write_data_reg;
   wire [3:0] reg_address;
   wire [7:0] read_data_reg;
   wire [7:0] reg0_A;
   wire [7:0] reg1_B;
   wire [7:0] reg2_config;
   wire [7:0] reg3_div_ratio;
   wire [3:0] alu_func;
   wire [15:0] alu_out;
   wire [7:0] rx_p_data;
   wire [7:0] data_to_fifo;
   wire [7:0] fifo_to_tx;
   wire [7:0] rx_out_data;
   wire [7:0] rx_div_ratio;
   wire SYNOPSYS_UNCONNECTED__0;
   wire SYNOPSYS_UNCONNECTED__1;
   wire SYNOPSYS_UNCONNECTED__2;
   wire SYNOPSYS_UNCONNECTED__3;

   assign SO[2] = rx_p_data[1] ;
   assign SO[0] = pulsing_empty ;

   // Module instantiations
   CLKINVX8M REF_CLK__L2_I0 (
	.Y(REF_CLK__L2_N0),
	.A(REF_CLK__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M REF_CLK__L1_I0 (
	.Y(REF_CLK__L1_N0),
	.A(REF_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX8M UART_CLK__L2_I0 (
	.Y(UART_CLK__L2_N0),
	.A(UART_CLK__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M UART_CLK__L1_I0 (
	.Y(UART_CLK__L1_N0),
	.A(UART_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX32M scan_clk__L12_I0 (
	.Y(scan_clk__L12_N0),
	.A(scan_clk__L11_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M scan_clk__L11_I0 (
	.Y(scan_clk__L11_N0),
	.A(scan_clk__L10_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX40M scan_clk__L10_I0 (
	.Y(scan_clk__L10_N0),
	.A(scan_clk__L9_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX40M scan_clk__L9_I1 (
	.Y(scan_clk__L9_N1),
	.A(scan_clk__L8_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX24M scan_clk__L9_I0 (
	.Y(scan_clk__L9_N0),
	.A(scan_clk__L8_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX40M scan_clk__L8_I1 (
	.Y(scan_clk__L8_N1),
	.A(scan_clk__L7_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX24M scan_clk__L8_I0 (
	.Y(scan_clk__L8_N0),
	.A(scan_clk__L7_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX40M scan_clk__L7_I1 (
	.Y(scan_clk__L7_N1),
	.A(scan_clk__L6_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX24M scan_clk__L7_I0 (
	.Y(scan_clk__L7_N0),
	.A(scan_clk__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX24M scan_clk__L6_I1 (
	.Y(scan_clk__L6_N1),
	.A(scan_clk__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX24M scan_clk__L6_I0 (
	.Y(scan_clk__L6_N0),
	.A(scan_clk__L5_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX24M scan_clk__L5_I1 (
	.Y(scan_clk__L5_N1),
	.A(scan_clk__L4_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX24M scan_clk__L5_I0 (
	.Y(scan_clk__L5_N0),
	.A(scan_clk__L4_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX24M scan_clk__L4_I0 (
	.Y(scan_clk__L4_N0),
	.A(scan_clk__L3_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX24M scan_clk__L3_I0 (
	.Y(scan_clk__L3_N0),
	.A(scan_clk__L2_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX16M scan_clk__L2_I0 (
	.Y(scan_clk__L2_N0),
	.A(scan_clk__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M scan_clk__L1_I0 (
	.Y(scan_clk__L1_N0),
	.A(scan_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M ref_clock__L5_I7 (
	.Y(ref_clock__L5_N7),
	.A(ref_clock__L4_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M ref_clock__L5_I6 (
	.Y(ref_clock__L5_N6),
	.A(ref_clock__L4_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M ref_clock__L5_I5 (
	.Y(ref_clock__L5_N5),
	.A(ref_clock__L4_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M ref_clock__L5_I4 (
	.Y(ref_clock__L5_N4),
	.A(ref_clock__L4_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M ref_clock__L5_I3 (
	.Y(ref_clock__L5_N3),
	.A(ref_clock__L4_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M ref_clock__L5_I2 (
	.Y(ref_clock__L5_N2),
	.A(ref_clock__L4_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M ref_clock__L5_I1 (
	.Y(ref_clock__L5_N1),
	.A(ref_clock__L4_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M ref_clock__L5_I0 (
	.Y(ref_clock__L5_N0),
	.A(ref_clock__L4_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M ref_clock__L4_I3 (
	.Y(ref_clock__L4_N3),
	.A(ref_clock__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M ref_clock__L4_I2 (
	.Y(ref_clock__L4_N2),
	.A(ref_clock__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M ref_clock__L4_I1 (
	.Y(ref_clock__L4_N1),
	.A(ref_clock__L3_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M ref_clock__L4_I0 (
	.Y(ref_clock__L4_N0),
	.A(ref_clock__L3_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M ref_clock__L3_I1 (
	.Y(ref_clock__L3_N1),
	.A(ref_clock__L2_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M ref_clock__L3_I0 (
	.Y(ref_clock__L3_N0),
	.A(ref_clock__L2_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M ref_clock__L2_I0 (
	.Y(ref_clock__L2_N0),
	.A(ref_clock__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX12M ref_clock__L1_I0 (
	.Y(ref_clock__L1_N0),
	.A(ref_clock), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX32M gated_clk__L3_I1 (
	.Y(gated_clk__L3_N1),
	.A(gated_clk__L2_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX32M gated_clk__L3_I0 (
	.Y(gated_clk__L3_N0),
	.A(gated_clk__L2_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX24M gated_clk__L2_I0 (
	.Y(gated_clk__L2_N0),
	.A(gated_clk__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX8M gated_clk__L1_I0 (
	.Y(gated_clk__L1_N0),
	.A(gated_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX24M uart_clock__L12_I1 (
	.Y(uart_clock__L12_N1),
	.A(uart_clock__L11_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX24M uart_clock__L12_I0 (
	.Y(uart_clock__L12_N0),
	.A(uart_clock__L11_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M uart_clock__L11_I0 (
	.Y(uart_clock__L11_N0),
	.A(uart_clock__L10_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M uart_clock__L10_I0 (
	.Y(uart_clock__L10_N0),
	.A(uart_clock__L9_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX40M uart_clock__L9_I0 (
	.Y(uart_clock__L9_N0),
	.A(uart_clock__L8_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M uart_clock__L8_I0 (
	.Y(uart_clock__L8_N0),
	.A(uart_clock__L7_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M uart_clock__L7_I2 (
	.Y(uart_clock__L7_N2),
	.A(uart_clock__L6_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX24M uart_clock__L7_I1 (
	.Y(uart_clock__L7_N1),
	.A(uart_clock__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX24M uart_clock__L7_I0 (
	.Y(uart_clock__L7_N0),
	.A(uart_clock__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M uart_clock__L6_I1 (
	.Y(uart_clock__L6_N1),
	.A(uart_clock__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M uart_clock__L6_I0 (
	.Y(uart_clock__L6_N0),
	.A(uart_clock__L5_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M uart_clock__L5_I1 (
	.Y(uart_clock__L5_N1),
	.A(uart_clock__L4_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX32M uart_clock__L5_I0 (
	.Y(uart_clock__L5_N0),
	.A(uart_clock__L4_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M uart_clock__L4_I0 (
	.Y(uart_clock__L4_N0),
	.A(uart_clock__L3_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M uart_clock__L3_I2 (
	.Y(uart_clock__L3_N2),
	.A(uart_clock__L2_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX24M uart_clock__L3_I1 (
	.Y(uart_clock__L3_N1),
	.A(uart_clock__L2_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX24M uart_clock__L3_I0 (
	.Y(uart_clock__L3_N0),
	.A(uart_clock__L2_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX32M uart_clock__L2_I0 (
	.Y(uart_clock__L2_N0),
	.A(uart_clock__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M uart_clock__L1_I0 (
	.Y(uart_clock__L1_N0),
	.A(uart_clock), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX8M n12__Exclude_0 (
	.Y(n12__Exclude_0_NET),
	.A(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX8M n11__Exclude_0 (
	.Y(n11__Exclude_0_NET),
	.A(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX24M tx_clock__L3_I3 (
	.Y(tx_clock__L3_N3),
	.A(tx_clock__L2_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX24M tx_clock__L3_I2 (
	.Y(tx_clock__L3_N2),
	.A(tx_clock__L2_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX24M tx_clock__L3_I1 (
	.Y(tx_clock__L3_N1),
	.A(tx_clock__L2_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX24M tx_clock__L3_I0 (
	.Y(tx_clock__L3_N0),
	.A(tx_clock__L2_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M tx_clock__L2_I0 (
	.Y(tx_clock__L2_N0),
	.A(tx_clock__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M tx_clock__L1_I0 (
	.Y(tx_clock__L1_N0),
	.A(tx_clock), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX24M rx_clock__L3_I3 (
	.Y(rx_clock__L3_N3),
	.A(rx_clock__L2_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX24M rx_clock__L3_I2 (
	.Y(rx_clock__L3_N2),
	.A(rx_clock__L2_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX24M rx_clock__L3_I1 (
	.Y(rx_clock__L3_N1),
	.A(rx_clock__L2_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX24M rx_clock__L3_I0 (
	.Y(rx_clock__L3_N0),
	.A(rx_clock__L2_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX32M rx_clock__L2_I0 (
	.Y(rx_clock__L2_N0),
	.A(rx_clock__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX12M rx_clock__L1_I0 (
	.Y(rx_clock__L1_N0),
	.A(rx_clock), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX4M FE_OFC5_SE (
	.Y(FE_OFN5_SE),
	.A(SE), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX4M FE_OFC2_rst_from_sync2 (
	.Y(FE_OFN2_rst_from_sync2),
	.A(rst_from_sync2), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX8M FE_OFC1_rst_from_sync1 (
	.Y(FE_OFN1_rst_from_sync1),
	.A(FE_OFN0_rst_from_sync1), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX10M FE_OFC0_rst_from_sync1 (
	.Y(FE_OFN0_rst_from_sync1),
	.A(rst_from_sync1), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U1 (
	.Y(n2),
	.A(reg_address[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX4M U2 (
	.Y(n3),
	.A(reg_address[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U7 (
	.Y(n1),
	.A(test_mode), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X4M U13 (
	.Y(n27),
	.A(n35), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X4M U14 (
	.Y(n28),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X4M U15 (
	.Y(n29),
	.A(n41), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U16 (
	.Y(n30),
	.A(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U17 (
	.Y(n31),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U18 (
	.Y(n32),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U19 (
	.Y(n33),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U20 (
	.Y(n34),
	.A(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U21 (
	.Y(n35),
	.A(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U22 (
	.Y(n36),
	.A(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U23 (
	.Y(n37),
	.A(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U24 (
	.Y(n38),
	.A(FE_OFN5_SE), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U25 (
	.Y(n39),
	.A(n38), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U26 (
	.Y(n40),
	.A(n38), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U27 (
	.Y(n41),
	.A(n38), 
	.VDD(VDD), 
	.VSS(VSS));
   mux2X1_1 refmux (
	.IN_0(REF_CLK__L2_N0),
	.IN_1(scan_clk__L9_N0),
	.SEL(n1),
	.OUT(ref_clock), 
	.VDD(VDD), 
	.VSS(VSS));
   mux2X1_5 uartmux (
	.IN_0(UART_CLK__L2_N0),
	.IN_1(scan_clk__L2_N0),
	.SEL(n1),
	.OUT(uart_clock), 
	.VDD(VDD), 
	.VSS(VSS));
   mux2X1_4 txmux (
	.IN_0(TX_CLK),
	.IN_1(scan_clk__L12_N0),
	.SEL(n1),
	.OUT(tx_clock), 
	.VDD(VDD), 
	.VSS(VSS));
   mux2X1_3 rxmux (
	.IN_0(RX_CLK),
	.IN_1(scan_clk__L12_N0),
	.SEL(n1),
	.OUT(rx_clock), 
	.VDD(VDD), 
	.VSS(VSS));
   mux2X1_2 rstmux (
	.IN_0(RST),
	.IN_1(scan_rst),
	.SEL(n1),
	.OUT(rst_to_sync), 
	.VDD(VDD), 
	.VSS(VSS));
   mux2X1_0 rst1mux (
	.IN_0(sync_rst1),
	.IN_1(scan_rst),
	.SEL(n1),
	.OUT(rst_from_sync1), 
	.VDD(VDD), 
	.VSS(VSS));
   mux2X1_6 rst2mux (
	.IN_0(sync_rst2),
	.IN_1(scan_rst),
	.SEL(n1),
	.OUT(rst_from_sync2), 
	.VDD(VDD), 
	.VSS(VSS));
   RegisterFile_test_1 RegFile (
	.WrData({ write_data_reg[7],
		write_data_reg[6],
		write_data_reg[5],
		write_data_reg[4],
		write_data_reg[3],
		write_data_reg[2],
		write_data_reg[1],
		write_data_reg[0] }),
	.Address({ reg_address[3],
		reg_address[2],
		n3,
		n2 }),
	.WrEn(write_enable_reg),
	.RdEn(read_enable_reg),
	.CLK(ref_clock__L5_N0),
	.RST(rst_from_sync1),
	.RdData({ read_data_reg[7],
		read_data_reg[6],
		read_data_reg[5],
		read_data_reg[4],
		read_data_reg[3],
		read_data_reg[2],
		read_data_reg[1],
		read_data_reg[0] }),
	.RdData_Valid(read_valid_reg),
	.REG0({ reg0_A[7],
		reg0_A[6],
		reg0_A[5],
		reg0_A[4],
		reg0_A[3],
		reg0_A[2],
		reg0_A[1],
		reg0_A[0] }),
	.REG1({ reg1_B[7],
		reg1_B[6],
		reg1_B[5],
		reg1_B[4],
		reg1_B[3],
		reg1_B[2],
		reg1_B[1],
		reg1_B[0] }),
	.REG2({ reg2_config[7],
		reg2_config[6],
		reg2_config[5],
		reg2_config[4],
		reg2_config[3],
		reg2_config[2],
		reg2_config[1],
		reg2_config[0] }),
	.REG3({ reg3_div_ratio[7],
		reg3_div_ratio[6],
		reg3_div_ratio[5],
		reg3_div_ratio[4],
		reg3_div_ratio[3],
		reg3_div_ratio[2],
		reg3_div_ratio[1],
		reg3_div_ratio[0] }),
	.test_si2(SI[2]),
	.test_si1(n25),
	.test_so2(n22),
	.test_so1(SO[3]),
	.test_se(FE_OFN5_SE),
	.FE_OFN0_rst_from_sync1(FE_OFN0_rst_from_sync1),
	.FE_OFN1_rst_from_sync1(FE_OFN1_rst_from_sync1),
	.ref_clock__L5_N4(ref_clock__L5_N4),
	.ref_clock__L5_N5(ref_clock__L5_N5),
	.ref_clock__L5_N6(ref_clock__L5_N6),
	.ref_clock__L5_N7(ref_clock__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   ALU_test_1 alu (
	.A({ reg0_A[7],
		reg0_A[6],
		reg0_A[5],
		reg0_A[4],
		reg0_A[3],
		reg0_A[2],
		reg0_A[1],
		reg0_A[0] }),
	.B({ reg1_B[7],
		reg1_B[6],
		reg1_B[5],
		reg1_B[4],
		reg1_B[3],
		reg1_B[2],
		reg1_B[1],
		reg1_B[0] }),
	.ALU_FUN({ alu_func[3],
		alu_func[2],
		alu_func[1],
		alu_func[0] }),
	.Enable(alu_enable),
	.CLK(gated_clk__L3_N0),
	.RST(FE_OFN1_rst_from_sync1),
	.ALU_OUT({ alu_out[15],
		alu_out[14],
		alu_out[13],
		alu_out[12],
		alu_out[11],
		alu_out[10],
		alu_out[9],
		alu_out[8],
		alu_out[7],
		alu_out[6],
		alu_out[5],
		alu_out[4],
		alu_out[3],
		alu_out[2],
		alu_out[1],
		alu_out[0] }),
	.OUT_VALID(out_valid),
	.test_si(n22),
	.test_se(n29),
	.gated_clk__L3_N1(gated_clk__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SYS_CTRL_test_1 FSM (
	.RX_D_VLD(rx_d_valid),
	.RX_P_Data({ rx_p_data[7],
		rx_p_data[6],
		rx_p_data[5],
		rx_p_data[4],
		rx_p_data[3],
		rx_p_data[2],
		rx_p_data[1],
		rx_p_data[0] }),
	.ALU_OUT({ alu_out[15],
		alu_out[14],
		alu_out[13],
		alu_out[12],
		alu_out[11],
		alu_out[10],
		alu_out[9],
		alu_out[8],
		alu_out[7],
		alu_out[6],
		alu_out[5],
		alu_out[4],
		alu_out[3],
		alu_out[2],
		alu_out[1],
		alu_out[0] }),
	.OUT_Valid(out_valid),
	.RdData({ read_data_reg[7],
		read_data_reg[6],
		read_data_reg[5],
		read_data_reg[4],
		read_data_reg[3],
		read_data_reg[2],
		read_data_reg[1],
		read_data_reg[0] }),
	.RdData_Valid(read_valid_reg),
	.CLK(ref_clock__L5_N0),
	.RST(rst_from_sync1),
	.fifo_full(full),
	.busyFall(tx_idle),
	.ALU_EN(alu_enable),
	.ALU_FUNC({ alu_func[3],
		alu_func[2],
		alu_func[1],
		alu_func[0] }),
	.CLK_EN(clock_gate_enable),
	.Address({ reg_address[3],
		reg_address[2],
		reg_address[1],
		reg_address[0] }),
	.WrEn(write_enable_reg),
	.RdEn(read_enable_reg),
	.WrData({ write_data_reg[7],
		write_data_reg[6],
		write_data_reg[5],
		write_data_reg[4],
		write_data_reg[3],
		write_data_reg[2],
		write_data_reg[1],
		write_data_reg[0] }),
	.TX_P_Data({ data_to_fifo[7],
		data_to_fifo[6],
		data_to_fifo[5],
		data_to_fifo[4],
		data_to_fifo[3],
		data_to_fifo[2],
		data_to_fifo[1],
		data_to_fifo[0] }),
	.TX_D_VLD(write_inc),
	.test_si(SI[3]),
	.test_so(n25),
	.test_se(n32),
	.FE_OFN1_rst_from_sync1(FE_OFN1_rst_from_sync1), 
	.VDD(VDD), 
	.VSS(VSS));
   FIFO_test_1 fifo (
	.W_CLK(ref_clock__L5_N1),
	.W_RST(rst_from_sync1),
	.W_INC(write_inc),
	.R_CLK(tx_clock__L3_N0),
	.R_RST(FE_OFN2_rst_from_sync2),
	.R_INC(read_inc),
	.WR_DATA({ data_to_fifo[7],
		data_to_fifo[6],
		data_to_fifo[5],
		data_to_fifo[4],
		data_to_fifo[3],
		data_to_fifo[2],
		data_to_fifo[1],
		data_to_fifo[0] }),
	.RD_DATA({ fifo_to_tx[7],
		fifo_to_tx[6],
		fifo_to_tx[5],
		fifo_to_tx[4],
		fifo_to_tx[3],
		fifo_to_tx[2],
		fifo_to_tx[1],
		fifo_to_tx[0] }),
	.full(full),
	.empty(empty),
	.test_si2(SI[0]),
	.test_si1(rx_p_data[7]),
	.test_so2(n17),
	.test_so1(SO[1]),
	.test_se(FE_OFN5_SE),
	.tx_clock__L3_N1(tx_clock__L3_N1),
	.tx_clock__L3_N2(tx_clock__L3_N2),
	.ref_clock__L5_N2(ref_clock__L5_N2),
	.ref_clock__L5_N3(ref_clock__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   UART_RX_test_1 rx (
	.RX_IN(RX_IN),
	.Prescale({ reg2_config[7],
		reg2_config[6],
		reg2_config[5],
		reg2_config[4],
		reg2_config[3],
		reg2_config[2] }),
	.PAR_EN(reg2_config[0]),
	.PAR_TYP(reg2_config[1]),
	.CLK(rx_clock__L3_N0),
	.RST(rst_from_sync2),
	.P_DATA({ rx_out_data[7],
		rx_out_data[6],
		rx_out_data[5],
		rx_out_data[4],
		rx_out_data[3],
		rx_out_data[2],
		rx_out_data[1],
		rx_out_data[0] }),
	.data_valid(rx_out_valid),
	.par_err(parity_error),
	.stp_err(frame_error),
	.test_si(n15),
	.test_so(n14),
	.test_se(n28),
	.rx_clock__L3_N1(rx_clock__L3_N1),
	.rx_clock__L3_N2(rx_clock__L3_N2),
	.rx_clock__L3_N3(rx_clock__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   UART_TX_test_1 tx (
	.clk(tx_clock__L3_N1),
	.rst(rst_from_sync2),
	.data({ fifo_to_tx[7],
		fifo_to_tx[6],
		fifo_to_tx[5],
		fifo_to_tx[4],
		fifo_to_tx[3],
		fifo_to_tx[2],
		fifo_to_tx[1],
		fifo_to_tx[0] }),
	.data_valid(vld),
	.parity_enable(reg2_config[0]),
	.parity_type(reg2_config[1]),
	.TX_OUT(TX_OUT),
	.busy(busy),
	.test_si(n14),
	.test_so(n13),
	.test_se(n27),
	.FE_OFN2_rst_from_sync2(FE_OFN2_rst_from_sync2),
	.tx_clock__L3_N2(tx_clock__L3_N2),
	.tx_clock__L3_N3(tx_clock__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DATA_SYNC_test_1 data_synch (
	.unsync_bus({ rx_out_data[7],
		rx_out_data[6],
		rx_out_data[5],
		rx_out_data[4],
		rx_out_data[3],
		rx_out_data[2],
		rx_out_data[1],
		rx_out_data[0] }),
	.bus_enable(rx_out_valid),
	.CLK(ref_clock__L5_N0),
	.RST(rst_from_sync1),
	.sync_bus({ rx_p_data[7],
		rx_p_data[6],
		rx_p_data[5],
		rx_p_data[4],
		rx_p_data[3],
		rx_p_data[2],
		rx_p_data[1],
		rx_p_data[0] }),
	.enable_pulse(rx_d_valid),
	.test_si2(SI[1]),
	.test_si1(n21),
	.test_se(n33),
	.ref_clock__L5_N1(ref_clock__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLK_GATE clkGate (
	.CLK_EN(clock_gate_enable),
	.CLK(ref_clock),
	.test_en(n1),
	.GATED_CLK(gated_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   PULSE_GEN_test_0 pulse_en (
	.CLK(tx_clock__L3_N1),
	.RST(FE_OFN2_rst_from_sync2),
	.LVL_SIG(busy),
	.PULSE_SIG(read_inc),
	.test_si(n17),
	.test_so(n16),
	.test_se(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   PULSE_GEN_test_1 pulse_valid (
	.CLK(tx_clock__L3_N1),
	.RST(FE_OFN2_rst_from_sync2),
	.LVL_SIG(pulsing_empty),
	.PULSE_SIG(vld),
	.test_si(n16),
	.test_so(n15),
	.test_se(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   PULSE_SAMEZERO_GEN_test_1 u7 (
	.CLK(tx_clock__L3_N0),
	.RST(FE_OFN2_rst_from_sync2),
	.busyFall(tx_idle),
	.empty(empty),
	.PULSE_SIG(pulsing_empty),
	.test_si(n9),
	.test_se(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   PULSE_NEG_GEN_test_1 busy_faling (
	.CLK(tx_clock__L3_N1),
	.RST(FE_OFN2_rst_from_sync2),
	.LVL_SIG(busy),
	.PULSE_SIG(tx_idle),
	.test_si(out_valid),
	.test_so(n21),
	.test_se(n36), 
	.VDD(VDD), 
	.VSS(VSS));
   ClkDiv_test_0 u0 (
	.i_ref_clk(uart_clock__L12_N1),
	.i_rst_n(rst_from_sync2),
	.i_clk_en(1'b1),
	.i_div_ratio({ reg3_div_ratio[7],
		reg3_div_ratio[6],
		reg3_div_ratio[5],
		reg3_div_ratio[4],
		reg3_div_ratio[3],
		reg3_div_ratio[2],
		reg3_div_ratio[1],
		reg3_div_ratio[0] }),
	.o_div_clk(TX_CLK),
	.test_si(n13),
	.test_so(n12),
	.test_se(n39),
	.n12__Exclude_0_NET(n12__Exclude_0_NET),
	.uart_clock__L3_N0(uart_clock__L3_N0),
	.uart_clock__L7_N0(uart_clock__L7_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   ClkDiv_test_1 u1 (
	.i_ref_clk(uart_clock__L12_N0),
	.i_rst_n(rst_from_sync2),
	.i_clk_en(1'b1),
	.i_div_ratio({ 1'b0,
		1'b0,
		1'b0,
		1'b0,
		rx_div_ratio[3],
		rx_div_ratio[2],
		rx_div_ratio[1],
		rx_div_ratio[0] }),
	.o_div_clk(RX_CLK),
	.test_si(n12__Exclude_0_NET),
	.test_so(n11),
	.test_se(n37),
	.n11__Exclude_0_NET(n11__Exclude_0_NET),
	.uart_clock__L3_N1(uart_clock__L3_N1),
	.uart_clock__L7_N1(uart_clock__L7_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   RST_SYNC_test_0 u2 (
	.CLK(ref_clock__L5_N1),
	.RST(rst_to_sync),
	.SYNC_RST(sync_rst1),
	.test_si(n11__Exclude_0_NET),
	.test_so(n10),
	.test_se(n36), 
	.VDD(VDD), 
	.VSS(VSS));
   RST_SYNC_test_1 u3 (
	.CLK(uart_clock__L12_N0),
	.RST(rst_to_sync),
	.SYNC_RST(sync_rst2),
	.test_si(n10),
	.test_so(n9),
	.test_se(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   custom_mux mux_prescale (
	.selector({ reg2_config[7],
		reg2_config[6],
		reg2_config[5],
		reg2_config[4],
		reg2_config[3],
		reg2_config[2] }),
	.div_ratio({ SYNOPSYS_UNCONNECTED__0,
		SYNOPSYS_UNCONNECTED__1,
		SYNOPSYS_UNCONNECTED__2,
		SYNOPSYS_UNCONNECTED__3,
		rx_div_ratio[3],
		rx_div_ratio[2],
		rx_div_ratio[1],
		rx_div_ratio[0] }), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

